-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     Jun 5 2019 04:46:17

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "latticehx1k" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of latticehx1k
entity latticehx1k is
port (
    led : out std_logic_vector(4 downto 0);
    o_serial_data : out std_logic;
    to_ir : out std_logic;
    sd : out std_logic;
    from_pc : in std_logic;
    clk_in : in std_logic);
end latticehx1k;

-- Architecture of latticehx1k
-- View name is \INTERFACE\
architecture \INTERFACE\ of latticehx1k is

signal \N__30236\ : std_logic;
signal \N__30235\ : std_logic;
signal \N__30234\ : std_logic;
signal \N__30227\ : std_logic;
signal \N__30226\ : std_logic;
signal \N__30225\ : std_logic;
signal \N__30218\ : std_logic;
signal \N__30217\ : std_logic;
signal \N__30216\ : std_logic;
signal \N__30209\ : std_logic;
signal \N__30208\ : std_logic;
signal \N__30207\ : std_logic;
signal \N__30200\ : std_logic;
signal \N__30199\ : std_logic;
signal \N__30198\ : std_logic;
signal \N__30191\ : std_logic;
signal \N__30190\ : std_logic;
signal \N__30189\ : std_logic;
signal \N__30182\ : std_logic;
signal \N__30181\ : std_logic;
signal \N__30180\ : std_logic;
signal \N__30173\ : std_logic;
signal \N__30172\ : std_logic;
signal \N__30171\ : std_logic;
signal \N__30164\ : std_logic;
signal \N__30163\ : std_logic;
signal \N__30162\ : std_logic;
signal \N__30155\ : std_logic;
signal \N__30154\ : std_logic;
signal \N__30153\ : std_logic;
signal \N__30136\ : std_logic;
signal \N__30133\ : std_logic;
signal \N__30130\ : std_logic;
signal \N__30127\ : std_logic;
signal \N__30124\ : std_logic;
signal \N__30121\ : std_logic;
signal \N__30120\ : std_logic;
signal \N__30119\ : std_logic;
signal \N__30118\ : std_logic;
signal \N__30113\ : std_logic;
signal \N__30108\ : std_logic;
signal \N__30107\ : std_logic;
signal \N__30104\ : std_logic;
signal \N__30101\ : std_logic;
signal \N__30098\ : std_logic;
signal \N__30095\ : std_logic;
signal \N__30092\ : std_logic;
signal \N__30089\ : std_logic;
signal \N__30082\ : std_logic;
signal \N__30081\ : std_logic;
signal \N__30078\ : std_logic;
signal \N__30075\ : std_logic;
signal \N__30074\ : std_logic;
signal \N__30073\ : std_logic;
signal \N__30072\ : std_logic;
signal \N__30069\ : std_logic;
signal \N__30066\ : std_logic;
signal \N__30061\ : std_logic;
signal \N__30058\ : std_logic;
signal \N__30055\ : std_logic;
signal \N__30046\ : std_logic;
signal \N__30043\ : std_logic;
signal \N__30040\ : std_logic;
signal \N__30039\ : std_logic;
signal \N__30038\ : std_logic;
signal \N__30037\ : std_logic;
signal \N__30034\ : std_logic;
signal \N__30031\ : std_logic;
signal \N__30030\ : std_logic;
signal \N__30029\ : std_logic;
signal \N__30028\ : std_logic;
signal \N__30027\ : std_logic;
signal \N__30024\ : std_logic;
signal \N__30021\ : std_logic;
signal \N__30016\ : std_logic;
signal \N__30013\ : std_logic;
signal \N__30006\ : std_logic;
signal \N__30003\ : std_logic;
signal \N__29992\ : std_logic;
signal \N__29989\ : std_logic;
signal \N__29988\ : std_logic;
signal \N__29987\ : std_logic;
signal \N__29986\ : std_logic;
signal \N__29985\ : std_logic;
signal \N__29982\ : std_logic;
signal \N__29977\ : std_logic;
signal \N__29972\ : std_logic;
signal \N__29969\ : std_logic;
signal \N__29962\ : std_logic;
signal \N__29961\ : std_logic;
signal \N__29960\ : std_logic;
signal \N__29959\ : std_logic;
signal \N__29958\ : std_logic;
signal \N__29957\ : std_logic;
signal \N__29956\ : std_logic;
signal \N__29953\ : std_logic;
signal \N__29952\ : std_logic;
signal \N__29951\ : std_logic;
signal \N__29950\ : std_logic;
signal \N__29945\ : std_logic;
signal \N__29940\ : std_logic;
signal \N__29939\ : std_logic;
signal \N__29936\ : std_logic;
signal \N__29929\ : std_logic;
signal \N__29924\ : std_logic;
signal \N__29921\ : std_logic;
signal \N__29918\ : std_logic;
signal \N__29915\ : std_logic;
signal \N__29912\ : std_logic;
signal \N__29905\ : std_logic;
signal \N__29902\ : std_logic;
signal \N__29893\ : std_logic;
signal \N__29892\ : std_logic;
signal \N__29891\ : std_logic;
signal \N__29888\ : std_logic;
signal \N__29883\ : std_logic;
signal \N__29882\ : std_logic;
signal \N__29877\ : std_logic;
signal \N__29874\ : std_logic;
signal \N__29869\ : std_logic;
signal \N__29868\ : std_logic;
signal \N__29867\ : std_logic;
signal \N__29864\ : std_logic;
signal \N__29859\ : std_logic;
signal \N__29854\ : std_logic;
signal \N__29851\ : std_logic;
signal \N__29848\ : std_logic;
signal \N__29845\ : std_logic;
signal \N__29844\ : std_logic;
signal \N__29843\ : std_logic;
signal \N__29840\ : std_logic;
signal \N__29837\ : std_logic;
signal \N__29832\ : std_logic;
signal \N__29829\ : std_logic;
signal \N__29826\ : std_logic;
signal \N__29821\ : std_logic;
signal \N__29820\ : std_logic;
signal \N__29817\ : std_logic;
signal \N__29816\ : std_logic;
signal \N__29815\ : std_logic;
signal \N__29814\ : std_logic;
signal \N__29813\ : std_logic;
signal \N__29812\ : std_logic;
signal \N__29809\ : std_logic;
signal \N__29806\ : std_logic;
signal \N__29799\ : std_logic;
signal \N__29794\ : std_logic;
signal \N__29791\ : std_logic;
signal \N__29782\ : std_logic;
signal \N__29781\ : std_logic;
signal \N__29780\ : std_logic;
signal \N__29779\ : std_logic;
signal \N__29778\ : std_logic;
signal \N__29775\ : std_logic;
signal \N__29774\ : std_logic;
signal \N__29773\ : std_logic;
signal \N__29768\ : std_logic;
signal \N__29765\ : std_logic;
signal \N__29762\ : std_logic;
signal \N__29761\ : std_logic;
signal \N__29758\ : std_logic;
signal \N__29755\ : std_logic;
signal \N__29752\ : std_logic;
signal \N__29749\ : std_logic;
signal \N__29744\ : std_logic;
signal \N__29741\ : std_logic;
signal \N__29736\ : std_logic;
signal \N__29733\ : std_logic;
signal \N__29726\ : std_logic;
signal \N__29725\ : std_logic;
signal \N__29724\ : std_logic;
signal \N__29721\ : std_logic;
signal \N__29718\ : std_logic;
signal \N__29715\ : std_logic;
signal \N__29710\ : std_logic;
signal \N__29701\ : std_logic;
signal \N__29700\ : std_logic;
signal \N__29699\ : std_logic;
signal \N__29696\ : std_logic;
signal \N__29693\ : std_logic;
signal \N__29690\ : std_logic;
signal \N__29689\ : std_logic;
signal \N__29686\ : std_logic;
signal \N__29685\ : std_logic;
signal \N__29684\ : std_logic;
signal \N__29683\ : std_logic;
signal \N__29678\ : std_logic;
signal \N__29675\ : std_logic;
signal \N__29672\ : std_logic;
signal \N__29665\ : std_logic;
signal \N__29660\ : std_logic;
signal \N__29653\ : std_logic;
signal \N__29650\ : std_logic;
signal \N__29647\ : std_logic;
signal \N__29644\ : std_logic;
signal \N__29641\ : std_logic;
signal \N__29638\ : std_logic;
signal \N__29637\ : std_logic;
signal \N__29634\ : std_logic;
signal \N__29631\ : std_logic;
signal \N__29630\ : std_logic;
signal \N__29629\ : std_logic;
signal \N__29624\ : std_logic;
signal \N__29619\ : std_logic;
signal \N__29616\ : std_logic;
signal \N__29613\ : std_logic;
signal \N__29612\ : std_logic;
signal \N__29609\ : std_logic;
signal \N__29606\ : std_logic;
signal \N__29603\ : std_logic;
signal \N__29596\ : std_logic;
signal \N__29593\ : std_logic;
signal \N__29590\ : std_logic;
signal \N__29587\ : std_logic;
signal \N__29584\ : std_logic;
signal \N__29581\ : std_logic;
signal \N__29578\ : std_logic;
signal \N__29577\ : std_logic;
signal \N__29576\ : std_logic;
signal \N__29575\ : std_logic;
signal \N__29574\ : std_logic;
signal \N__29573\ : std_logic;
signal \N__29572\ : std_logic;
signal \N__29569\ : std_logic;
signal \N__29562\ : std_logic;
signal \N__29555\ : std_logic;
signal \N__29548\ : std_logic;
signal \N__29547\ : std_logic;
signal \N__29546\ : std_logic;
signal \N__29541\ : std_logic;
signal \N__29540\ : std_logic;
signal \N__29539\ : std_logic;
signal \N__29536\ : std_logic;
signal \N__29533\ : std_logic;
signal \N__29532\ : std_logic;
signal \N__29529\ : std_logic;
signal \N__29526\ : std_logic;
signal \N__29521\ : std_logic;
signal \N__29518\ : std_logic;
signal \N__29513\ : std_logic;
signal \N__29512\ : std_logic;
signal \N__29509\ : std_logic;
signal \N__29506\ : std_logic;
signal \N__29503\ : std_logic;
signal \N__29500\ : std_logic;
signal \N__29491\ : std_logic;
signal \N__29490\ : std_logic;
signal \N__29487\ : std_logic;
signal \N__29484\ : std_logic;
signal \N__29481\ : std_logic;
signal \N__29480\ : std_logic;
signal \N__29479\ : std_logic;
signal \N__29478\ : std_logic;
signal \N__29477\ : std_logic;
signal \N__29476\ : std_logic;
signal \N__29475\ : std_logic;
signal \N__29474\ : std_logic;
signal \N__29473\ : std_logic;
signal \N__29472\ : std_logic;
signal \N__29471\ : std_logic;
signal \N__29470\ : std_logic;
signal \N__29469\ : std_logic;
signal \N__29468\ : std_logic;
signal \N__29467\ : std_logic;
signal \N__29466\ : std_logic;
signal \N__29465\ : std_logic;
signal \N__29464\ : std_logic;
signal \N__29463\ : std_logic;
signal \N__29462\ : std_logic;
signal \N__29461\ : std_logic;
signal \N__29460\ : std_logic;
signal \N__29459\ : std_logic;
signal \N__29458\ : std_logic;
signal \N__29457\ : std_logic;
signal \N__29456\ : std_logic;
signal \N__29455\ : std_logic;
signal \N__29454\ : std_logic;
signal \N__29453\ : std_logic;
signal \N__29452\ : std_logic;
signal \N__29451\ : std_logic;
signal \N__29450\ : std_logic;
signal \N__29449\ : std_logic;
signal \N__29448\ : std_logic;
signal \N__29447\ : std_logic;
signal \N__29446\ : std_logic;
signal \N__29445\ : std_logic;
signal \N__29444\ : std_logic;
signal \N__29443\ : std_logic;
signal \N__29442\ : std_logic;
signal \N__29441\ : std_logic;
signal \N__29440\ : std_logic;
signal \N__29439\ : std_logic;
signal \N__29438\ : std_logic;
signal \N__29437\ : std_logic;
signal \N__29436\ : std_logic;
signal \N__29435\ : std_logic;
signal \N__29434\ : std_logic;
signal \N__29433\ : std_logic;
signal \N__29432\ : std_logic;
signal \N__29431\ : std_logic;
signal \N__29430\ : std_logic;
signal \N__29429\ : std_logic;
signal \N__29428\ : std_logic;
signal \N__29427\ : std_logic;
signal \N__29426\ : std_logic;
signal \N__29425\ : std_logic;
signal \N__29424\ : std_logic;
signal \N__29423\ : std_logic;
signal \N__29422\ : std_logic;
signal \N__29421\ : std_logic;
signal \N__29420\ : std_logic;
signal \N__29419\ : std_logic;
signal \N__29418\ : std_logic;
signal \N__29417\ : std_logic;
signal \N__29416\ : std_logic;
signal \N__29415\ : std_logic;
signal \N__29414\ : std_logic;
signal \N__29413\ : std_logic;
signal \N__29412\ : std_logic;
signal \N__29411\ : std_logic;
signal \N__29410\ : std_logic;
signal \N__29409\ : std_logic;
signal \N__29408\ : std_logic;
signal \N__29407\ : std_logic;
signal \N__29406\ : std_logic;
signal \N__29405\ : std_logic;
signal \N__29404\ : std_logic;
signal \N__29403\ : std_logic;
signal \N__29402\ : std_logic;
signal \N__29401\ : std_logic;
signal \N__29400\ : std_logic;
signal \N__29399\ : std_logic;
signal \N__29398\ : std_logic;
signal \N__29397\ : std_logic;
signal \N__29396\ : std_logic;
signal \N__29395\ : std_logic;
signal \N__29394\ : std_logic;
signal \N__29393\ : std_logic;
signal \N__29392\ : std_logic;
signal \N__29391\ : std_logic;
signal \N__29390\ : std_logic;
signal \N__29389\ : std_logic;
signal \N__29388\ : std_logic;
signal \N__29387\ : std_logic;
signal \N__29386\ : std_logic;
signal \N__29385\ : std_logic;
signal \N__29384\ : std_logic;
signal \N__29383\ : std_logic;
signal \N__29382\ : std_logic;
signal \N__29381\ : std_logic;
signal \N__29380\ : std_logic;
signal \N__29379\ : std_logic;
signal \N__29378\ : std_logic;
signal \N__29377\ : std_logic;
signal \N__29376\ : std_logic;
signal \N__29375\ : std_logic;
signal \N__29374\ : std_logic;
signal \N__29373\ : std_logic;
signal \N__29372\ : std_logic;
signal \N__29371\ : std_logic;
signal \N__29370\ : std_logic;
signal \N__29367\ : std_logic;
signal \N__29364\ : std_logic;
signal \N__29137\ : std_logic;
signal \N__29134\ : std_logic;
signal \N__29131\ : std_logic;
signal \N__29130\ : std_logic;
signal \N__29127\ : std_logic;
signal \N__29126\ : std_logic;
signal \N__29123\ : std_logic;
signal \N__29120\ : std_logic;
signal \N__29115\ : std_logic;
signal \N__29110\ : std_logic;
signal \N__29107\ : std_logic;
signal \N__29106\ : std_logic;
signal \N__29105\ : std_logic;
signal \N__29104\ : std_logic;
signal \N__29103\ : std_logic;
signal \N__29102\ : std_logic;
signal \N__29099\ : std_logic;
signal \N__29098\ : std_logic;
signal \N__29097\ : std_logic;
signal \N__29094\ : std_logic;
signal \N__29091\ : std_logic;
signal \N__29086\ : std_logic;
signal \N__29083\ : std_logic;
signal \N__29080\ : std_logic;
signal \N__29077\ : std_logic;
signal \N__29074\ : std_logic;
signal \N__29073\ : std_logic;
signal \N__29070\ : std_logic;
signal \N__29065\ : std_logic;
signal \N__29064\ : std_logic;
signal \N__29063\ : std_logic;
signal \N__29062\ : std_logic;
signal \N__29059\ : std_logic;
signal \N__29052\ : std_logic;
signal \N__29049\ : std_logic;
signal \N__29048\ : std_logic;
signal \N__29047\ : std_logic;
signal \N__29042\ : std_logic;
signal \N__29035\ : std_logic;
signal \N__29030\ : std_logic;
signal \N__29027\ : std_logic;
signal \N__29026\ : std_logic;
signal \N__29023\ : std_logic;
signal \N__29020\ : std_logic;
signal \N__29015\ : std_logic;
signal \N__29010\ : std_logic;
signal \N__29003\ : std_logic;
signal \N__28996\ : std_logic;
signal \N__28995\ : std_logic;
signal \N__28994\ : std_logic;
signal \N__28991\ : std_logic;
signal \N__28988\ : std_logic;
signal \N__28987\ : std_logic;
signal \N__28986\ : std_logic;
signal \N__28985\ : std_logic;
signal \N__28984\ : std_logic;
signal \N__28983\ : std_logic;
signal \N__28982\ : std_logic;
signal \N__28981\ : std_logic;
signal \N__28980\ : std_logic;
signal \N__28979\ : std_logic;
signal \N__28978\ : std_logic;
signal \N__28975\ : std_logic;
signal \N__28974\ : std_logic;
signal \N__28971\ : std_logic;
signal \N__28968\ : std_logic;
signal \N__28965\ : std_logic;
signal \N__28964\ : std_logic;
signal \N__28957\ : std_logic;
signal \N__28954\ : std_logic;
signal \N__28951\ : std_logic;
signal \N__28948\ : std_logic;
signal \N__28947\ : std_logic;
signal \N__28944\ : std_logic;
signal \N__28943\ : std_logic;
signal \N__28938\ : std_logic;
signal \N__28935\ : std_logic;
signal \N__28932\ : std_logic;
signal \N__28925\ : std_logic;
signal \N__28924\ : std_logic;
signal \N__28921\ : std_logic;
signal \N__28916\ : std_logic;
signal \N__28913\ : std_logic;
signal \N__28910\ : std_logic;
signal \N__28907\ : std_logic;
signal \N__28906\ : std_logic;
signal \N__28905\ : std_logic;
signal \N__28902\ : std_logic;
signal \N__28899\ : std_logic;
signal \N__28896\ : std_logic;
signal \N__28893\ : std_logic;
signal \N__28890\ : std_logic;
signal \N__28887\ : std_logic;
signal \N__28884\ : std_logic;
signal \N__28881\ : std_logic;
signal \N__28878\ : std_logic;
signal \N__28873\ : std_logic;
signal \N__28870\ : std_logic;
signal \N__28867\ : std_logic;
signal \N__28864\ : std_logic;
signal \N__28861\ : std_logic;
signal \N__28858\ : std_logic;
signal \N__28851\ : std_logic;
signal \N__28844\ : std_logic;
signal \N__28837\ : std_logic;
signal \N__28822\ : std_logic;
signal \N__28821\ : std_logic;
signal \N__28820\ : std_logic;
signal \N__28819\ : std_logic;
signal \N__28818\ : std_logic;
signal \N__28817\ : std_logic;
signal \N__28816\ : std_logic;
signal \N__28813\ : std_logic;
signal \N__28812\ : std_logic;
signal \N__28809\ : std_logic;
signal \N__28806\ : std_logic;
signal \N__28803\ : std_logic;
signal \N__28800\ : std_logic;
signal \N__28797\ : std_logic;
signal \N__28796\ : std_logic;
signal \N__28795\ : std_logic;
signal \N__28792\ : std_logic;
signal \N__28789\ : std_logic;
signal \N__28786\ : std_logic;
signal \N__28783\ : std_logic;
signal \N__28776\ : std_logic;
signal \N__28773\ : std_logic;
signal \N__28772\ : std_logic;
signal \N__28771\ : std_logic;
signal \N__28766\ : std_logic;
signal \N__28763\ : std_logic;
signal \N__28760\ : std_logic;
signal \N__28757\ : std_logic;
signal \N__28756\ : std_logic;
signal \N__28755\ : std_logic;
signal \N__28754\ : std_logic;
signal \N__28753\ : std_logic;
signal \N__28750\ : std_logic;
signal \N__28747\ : std_logic;
signal \N__28744\ : std_logic;
signal \N__28743\ : std_logic;
signal \N__28738\ : std_logic;
signal \N__28735\ : std_logic;
signal \N__28732\ : std_logic;
signal \N__28729\ : std_logic;
signal \N__28726\ : std_logic;
signal \N__28721\ : std_logic;
signal \N__28718\ : std_logic;
signal \N__28715\ : std_logic;
signal \N__28708\ : std_logic;
signal \N__28705\ : std_logic;
signal \N__28684\ : std_logic;
signal \N__28683\ : std_logic;
signal \N__28682\ : std_logic;
signal \N__28679\ : std_logic;
signal \N__28678\ : std_logic;
signal \N__28677\ : std_logic;
signal \N__28672\ : std_logic;
signal \N__28669\ : std_logic;
signal \N__28666\ : std_logic;
signal \N__28665\ : std_logic;
signal \N__28664\ : std_logic;
signal \N__28661\ : std_logic;
signal \N__28660\ : std_logic;
signal \N__28653\ : std_logic;
signal \N__28644\ : std_logic;
signal \N__28641\ : std_logic;
signal \N__28636\ : std_logic;
signal \N__28635\ : std_logic;
signal \N__28634\ : std_logic;
signal \N__28633\ : std_logic;
signal \N__28624\ : std_logic;
signal \N__28621\ : std_logic;
signal \N__28618\ : std_logic;
signal \N__28615\ : std_logic;
signal \N__28614\ : std_logic;
signal \N__28613\ : std_logic;
signal \N__28612\ : std_logic;
signal \N__28611\ : std_logic;
signal \N__28610\ : std_logic;
signal \N__28609\ : std_logic;
signal \N__28608\ : std_logic;
signal \N__28607\ : std_logic;
signal \N__28606\ : std_logic;
signal \N__28603\ : std_logic;
signal \N__28602\ : std_logic;
signal \N__28601\ : std_logic;
signal \N__28598\ : std_logic;
signal \N__28597\ : std_logic;
signal \N__28596\ : std_logic;
signal \N__28593\ : std_logic;
signal \N__28590\ : std_logic;
signal \N__28585\ : std_logic;
signal \N__28580\ : std_logic;
signal \N__28577\ : std_logic;
signal \N__28574\ : std_logic;
signal \N__28573\ : std_logic;
signal \N__28570\ : std_logic;
signal \N__28567\ : std_logic;
signal \N__28564\ : std_logic;
signal \N__28563\ : std_logic;
signal \N__28560\ : std_logic;
signal \N__28557\ : std_logic;
signal \N__28554\ : std_logic;
signal \N__28551\ : std_logic;
signal \N__28548\ : std_logic;
signal \N__28543\ : std_logic;
signal \N__28540\ : std_logic;
signal \N__28539\ : std_logic;
signal \N__28536\ : std_logic;
signal \N__28533\ : std_logic;
signal \N__28530\ : std_logic;
signal \N__28527\ : std_logic;
signal \N__28524\ : std_logic;
signal \N__28521\ : std_logic;
signal \N__28518\ : std_logic;
signal \N__28515\ : std_logic;
signal \N__28510\ : std_logic;
signal \N__28509\ : std_logic;
signal \N__28508\ : std_logic;
signal \N__28507\ : std_logic;
signal \N__28500\ : std_logic;
signal \N__28497\ : std_logic;
signal \N__28494\ : std_logic;
signal \N__28485\ : std_logic;
signal \N__28476\ : std_logic;
signal \N__28469\ : std_logic;
signal \N__28456\ : std_logic;
signal \N__28455\ : std_logic;
signal \N__28452\ : std_logic;
signal \N__28449\ : std_logic;
signal \N__28448\ : std_logic;
signal \N__28447\ : std_logic;
signal \N__28446\ : std_logic;
signal \N__28443\ : std_logic;
signal \N__28440\ : std_logic;
signal \N__28437\ : std_logic;
signal \N__28436\ : std_logic;
signal \N__28433\ : std_logic;
signal \N__28430\ : std_logic;
signal \N__28423\ : std_logic;
signal \N__28420\ : std_logic;
signal \N__28419\ : std_logic;
signal \N__28416\ : std_logic;
signal \N__28413\ : std_logic;
signal \N__28408\ : std_logic;
signal \N__28405\ : std_logic;
signal \N__28402\ : std_logic;
signal \N__28399\ : std_logic;
signal \N__28396\ : std_logic;
signal \N__28393\ : std_logic;
signal \N__28390\ : std_logic;
signal \N__28387\ : std_logic;
signal \N__28384\ : std_logic;
signal \N__28381\ : std_logic;
signal \N__28378\ : std_logic;
signal \N__28375\ : std_logic;
signal \N__28372\ : std_logic;
signal \N__28369\ : std_logic;
signal \N__28360\ : std_logic;
signal \N__28357\ : std_logic;
signal \N__28356\ : std_logic;
signal \N__28355\ : std_logic;
signal \N__28354\ : std_logic;
signal \N__28353\ : std_logic;
signal \N__28350\ : std_logic;
signal \N__28347\ : std_logic;
signal \N__28344\ : std_logic;
signal \N__28341\ : std_logic;
signal \N__28336\ : std_logic;
signal \N__28333\ : std_logic;
signal \N__28330\ : std_logic;
signal \N__28327\ : std_logic;
signal \N__28324\ : std_logic;
signal \N__28321\ : std_logic;
signal \N__28318\ : std_logic;
signal \N__28315\ : std_logic;
signal \N__28312\ : std_logic;
signal \N__28309\ : std_logic;
signal \N__28304\ : std_logic;
signal \N__28297\ : std_logic;
signal \N__28296\ : std_logic;
signal \N__28295\ : std_logic;
signal \N__28290\ : std_logic;
signal \N__28287\ : std_logic;
signal \N__28286\ : std_logic;
signal \N__28285\ : std_logic;
signal \N__28282\ : std_logic;
signal \N__28279\ : std_logic;
signal \N__28274\ : std_logic;
signal \N__28271\ : std_logic;
signal \N__28264\ : std_logic;
signal \N__28261\ : std_logic;
signal \N__28258\ : std_logic;
signal \N__28255\ : std_logic;
signal \N__28252\ : std_logic;
signal \N__28251\ : std_logic;
signal \N__28248\ : std_logic;
signal \N__28247\ : std_logic;
signal \N__28244\ : std_logic;
signal \N__28241\ : std_logic;
signal \N__28240\ : std_logic;
signal \N__28237\ : std_logic;
signal \N__28234\ : std_logic;
signal \N__28231\ : std_logic;
signal \N__28228\ : std_logic;
signal \N__28225\ : std_logic;
signal \N__28222\ : std_logic;
signal \N__28213\ : std_logic;
signal \N__28210\ : std_logic;
signal \N__28207\ : std_logic;
signal \N__28204\ : std_logic;
signal \N__28201\ : std_logic;
signal \N__28198\ : std_logic;
signal \N__28197\ : std_logic;
signal \N__28196\ : std_logic;
signal \N__28193\ : std_logic;
signal \N__28188\ : std_logic;
signal \N__28185\ : std_logic;
signal \N__28180\ : std_logic;
signal \N__28179\ : std_logic;
signal \N__28176\ : std_logic;
signal \N__28175\ : std_logic;
signal \N__28174\ : std_logic;
signal \N__28173\ : std_logic;
signal \N__28172\ : std_logic;
signal \N__28171\ : std_logic;
signal \N__28168\ : std_logic;
signal \N__28165\ : std_logic;
signal \N__28162\ : std_logic;
signal \N__28161\ : std_logic;
signal \N__28156\ : std_logic;
signal \N__28151\ : std_logic;
signal \N__28148\ : std_logic;
signal \N__28145\ : std_logic;
signal \N__28140\ : std_logic;
signal \N__28129\ : std_logic;
signal \N__28126\ : std_logic;
signal \N__28125\ : std_logic;
signal \N__28124\ : std_logic;
signal \N__28123\ : std_logic;
signal \N__28120\ : std_logic;
signal \N__28117\ : std_logic;
signal \N__28112\ : std_logic;
signal \N__28105\ : std_logic;
signal \N__28104\ : std_logic;
signal \N__28103\ : std_logic;
signal \N__28102\ : std_logic;
signal \N__28099\ : std_logic;
signal \N__28096\ : std_logic;
signal \N__28093\ : std_logic;
signal \N__28092\ : std_logic;
signal \N__28089\ : std_logic;
signal \N__28088\ : std_logic;
signal \N__28085\ : std_logic;
signal \N__28082\ : std_logic;
signal \N__28077\ : std_logic;
signal \N__28072\ : std_logic;
signal \N__28067\ : std_logic;
signal \N__28060\ : std_logic;
signal \N__28059\ : std_logic;
signal \N__28056\ : std_logic;
signal \N__28055\ : std_logic;
signal \N__28052\ : std_logic;
signal \N__28051\ : std_logic;
signal \N__28050\ : std_logic;
signal \N__28049\ : std_logic;
signal \N__28040\ : std_logic;
signal \N__28035\ : std_logic;
signal \N__28030\ : std_logic;
signal \N__28027\ : std_logic;
signal \N__28024\ : std_logic;
signal \N__28023\ : std_logic;
signal \N__28022\ : std_logic;
signal \N__28021\ : std_logic;
signal \N__28020\ : std_logic;
signal \N__28019\ : std_logic;
signal \N__28016\ : std_logic;
signal \N__28013\ : std_logic;
signal \N__28010\ : std_logic;
signal \N__28007\ : std_logic;
signal \N__28002\ : std_logic;
signal \N__27999\ : std_logic;
signal \N__27996\ : std_logic;
signal \N__27991\ : std_logic;
signal \N__27982\ : std_logic;
signal \N__27981\ : std_logic;
signal \N__27980\ : std_logic;
signal \N__27979\ : std_logic;
signal \N__27972\ : std_logic;
signal \N__27969\ : std_logic;
signal \N__27964\ : std_logic;
signal \N__27961\ : std_logic;
signal \N__27958\ : std_logic;
signal \N__27955\ : std_logic;
signal \N__27952\ : std_logic;
signal \N__27949\ : std_logic;
signal \N__27948\ : std_logic;
signal \N__27947\ : std_logic;
signal \N__27944\ : std_logic;
signal \N__27943\ : std_logic;
signal \N__27942\ : std_logic;
signal \N__27939\ : std_logic;
signal \N__27938\ : std_logic;
signal \N__27935\ : std_logic;
signal \N__27934\ : std_logic;
signal \N__27931\ : std_logic;
signal \N__27926\ : std_logic;
signal \N__27923\ : std_logic;
signal \N__27920\ : std_logic;
signal \N__27917\ : std_logic;
signal \N__27914\ : std_logic;
signal \N__27911\ : std_logic;
signal \N__27908\ : std_logic;
signal \N__27905\ : std_logic;
signal \N__27892\ : std_logic;
signal \N__27889\ : std_logic;
signal \N__27886\ : std_logic;
signal \N__27883\ : std_logic;
signal \N__27880\ : std_logic;
signal \N__27877\ : std_logic;
signal \N__27874\ : std_logic;
signal \N__27873\ : std_logic;
signal \N__27872\ : std_logic;
signal \N__27871\ : std_logic;
signal \N__27870\ : std_logic;
signal \N__27869\ : std_logic;
signal \N__27864\ : std_logic;
signal \N__27861\ : std_logic;
signal \N__27858\ : std_logic;
signal \N__27855\ : std_logic;
signal \N__27852\ : std_logic;
signal \N__27847\ : std_logic;
signal \N__27842\ : std_logic;
signal \N__27837\ : std_logic;
signal \N__27832\ : std_logic;
signal \N__27829\ : std_logic;
signal \N__27826\ : std_logic;
signal \N__27823\ : std_logic;
signal \N__27820\ : std_logic;
signal \N__27817\ : std_logic;
signal \N__27814\ : std_logic;
signal \N__27813\ : std_logic;
signal \N__27812\ : std_logic;
signal \N__27811\ : std_logic;
signal \N__27810\ : std_logic;
signal \N__27809\ : std_logic;
signal \N__27808\ : std_logic;
signal \N__27807\ : std_logic;
signal \N__27806\ : std_logic;
signal \N__27803\ : std_logic;
signal \N__27802\ : std_logic;
signal \N__27799\ : std_logic;
signal \N__27796\ : std_logic;
signal \N__27795\ : std_logic;
signal \N__27794\ : std_logic;
signal \N__27793\ : std_logic;
signal \N__27792\ : std_logic;
signal \N__27791\ : std_logic;
signal \N__27790\ : std_logic;
signal \N__27789\ : std_logic;
signal \N__27788\ : std_logic;
signal \N__27787\ : std_logic;
signal \N__27784\ : std_logic;
signal \N__27783\ : std_logic;
signal \N__27782\ : std_logic;
signal \N__27781\ : std_logic;
signal \N__27778\ : std_logic;
signal \N__27777\ : std_logic;
signal \N__27774\ : std_logic;
signal \N__27773\ : std_logic;
signal \N__27766\ : std_logic;
signal \N__27761\ : std_logic;
signal \N__27756\ : std_logic;
signal \N__27749\ : std_logic;
signal \N__27748\ : std_logic;
signal \N__27747\ : std_logic;
signal \N__27746\ : std_logic;
signal \N__27745\ : std_logic;
signal \N__27740\ : std_logic;
signal \N__27735\ : std_logic;
signal \N__27732\ : std_logic;
signal \N__27731\ : std_logic;
signal \N__27730\ : std_logic;
signal \N__27729\ : std_logic;
signal \N__27726\ : std_logic;
signal \N__27725\ : std_logic;
signal \N__27722\ : std_logic;
signal \N__27717\ : std_logic;
signal \N__27716\ : std_logic;
signal \N__27713\ : std_logic;
signal \N__27712\ : std_logic;
signal \N__27711\ : std_logic;
signal \N__27710\ : std_logic;
signal \N__27705\ : std_logic;
signal \N__27702\ : std_logic;
signal \N__27701\ : std_logic;
signal \N__27700\ : std_logic;
signal \N__27697\ : std_logic;
signal \N__27692\ : std_logic;
signal \N__27687\ : std_logic;
signal \N__27684\ : std_logic;
signal \N__27677\ : std_logic;
signal \N__27672\ : std_logic;
signal \N__27665\ : std_logic;
signal \N__27662\ : std_logic;
signal \N__27659\ : std_logic;
signal \N__27656\ : std_logic;
signal \N__27651\ : std_logic;
signal \N__27648\ : std_logic;
signal \N__27647\ : std_logic;
signal \N__27646\ : std_logic;
signal \N__27645\ : std_logic;
signal \N__27644\ : std_logic;
signal \N__27643\ : std_logic;
signal \N__27640\ : std_logic;
signal \N__27637\ : std_logic;
signal \N__27632\ : std_logic;
signal \N__27629\ : std_logic;
signal \N__27626\ : std_logic;
signal \N__27621\ : std_logic;
signal \N__27612\ : std_logic;
signal \N__27605\ : std_logic;
signal \N__27594\ : std_logic;
signal \N__27583\ : std_logic;
signal \N__27562\ : std_logic;
signal \N__27561\ : std_logic;
signal \N__27560\ : std_logic;
signal \N__27559\ : std_logic;
signal \N__27556\ : std_logic;
signal \N__27553\ : std_logic;
signal \N__27552\ : std_logic;
signal \N__27551\ : std_logic;
signal \N__27546\ : std_logic;
signal \N__27545\ : std_logic;
signal \N__27544\ : std_logic;
signal \N__27543\ : std_logic;
signal \N__27542\ : std_logic;
signal \N__27541\ : std_logic;
signal \N__27538\ : std_logic;
signal \N__27535\ : std_logic;
signal \N__27532\ : std_logic;
signal \N__27529\ : std_logic;
signal \N__27526\ : std_logic;
signal \N__27521\ : std_logic;
signal \N__27518\ : std_logic;
signal \N__27517\ : std_logic;
signal \N__27512\ : std_logic;
signal \N__27511\ : std_logic;
signal \N__27510\ : std_logic;
signal \N__27507\ : std_logic;
signal \N__27504\ : std_logic;
signal \N__27501\ : std_logic;
signal \N__27498\ : std_logic;
signal \N__27493\ : std_logic;
signal \N__27490\ : std_logic;
signal \N__27487\ : std_logic;
signal \N__27484\ : std_logic;
signal \N__27483\ : std_logic;
signal \N__27482\ : std_logic;
signal \N__27479\ : std_logic;
signal \N__27476\ : std_logic;
signal \N__27475\ : std_logic;
signal \N__27468\ : std_logic;
signal \N__27461\ : std_logic;
signal \N__27456\ : std_logic;
signal \N__27445\ : std_logic;
signal \N__27436\ : std_logic;
signal \N__27435\ : std_logic;
signal \N__27430\ : std_logic;
signal \N__27427\ : std_logic;
signal \N__27424\ : std_logic;
signal \N__27421\ : std_logic;
signal \N__27418\ : std_logic;
signal \N__27415\ : std_logic;
signal \N__27414\ : std_logic;
signal \N__27413\ : std_logic;
signal \N__27408\ : std_logic;
signal \N__27405\ : std_logic;
signal \N__27402\ : std_logic;
signal \N__27399\ : std_logic;
signal \N__27396\ : std_logic;
signal \N__27395\ : std_logic;
signal \N__27392\ : std_logic;
signal \N__27389\ : std_logic;
signal \N__27388\ : std_logic;
signal \N__27385\ : std_logic;
signal \N__27382\ : std_logic;
signal \N__27379\ : std_logic;
signal \N__27374\ : std_logic;
signal \N__27367\ : std_logic;
signal \N__27364\ : std_logic;
signal \N__27361\ : std_logic;
signal \N__27358\ : std_logic;
signal \N__27355\ : std_logic;
signal \N__27354\ : std_logic;
signal \N__27353\ : std_logic;
signal \N__27346\ : std_logic;
signal \N__27345\ : std_logic;
signal \N__27342\ : std_logic;
signal \N__27341\ : std_logic;
signal \N__27338\ : std_logic;
signal \N__27335\ : std_logic;
signal \N__27332\ : std_logic;
signal \N__27325\ : std_logic;
signal \N__27324\ : std_logic;
signal \N__27321\ : std_logic;
signal \N__27316\ : std_logic;
signal \N__27313\ : std_logic;
signal \N__27310\ : std_logic;
signal \N__27307\ : std_logic;
signal \N__27304\ : std_logic;
signal \N__27301\ : std_logic;
signal \N__27300\ : std_logic;
signal \N__27299\ : std_logic;
signal \N__27298\ : std_logic;
signal \N__27297\ : std_logic;
signal \N__27296\ : std_logic;
signal \N__27295\ : std_logic;
signal \N__27294\ : std_logic;
signal \N__27293\ : std_logic;
signal \N__27292\ : std_logic;
signal \N__27289\ : std_logic;
signal \N__27286\ : std_logic;
signal \N__27285\ : std_logic;
signal \N__27284\ : std_logic;
signal \N__27281\ : std_logic;
signal \N__27278\ : std_logic;
signal \N__27277\ : std_logic;
signal \N__27276\ : std_logic;
signal \N__27271\ : std_logic;
signal \N__27264\ : std_logic;
signal \N__27261\ : std_logic;
signal \N__27258\ : std_logic;
signal \N__27255\ : std_logic;
signal \N__27250\ : std_logic;
signal \N__27249\ : std_logic;
signal \N__27248\ : std_logic;
signal \N__27247\ : std_logic;
signal \N__27246\ : std_logic;
signal \N__27243\ : std_logic;
signal \N__27240\ : std_logic;
signal \N__27235\ : std_logic;
signal \N__27232\ : std_logic;
signal \N__27227\ : std_logic;
signal \N__27220\ : std_logic;
signal \N__27213\ : std_logic;
signal \N__27212\ : std_logic;
signal \N__27211\ : std_logic;
signal \N__27210\ : std_logic;
signal \N__27209\ : std_logic;
signal \N__27206\ : std_logic;
signal \N__27201\ : std_logic;
signal \N__27194\ : std_logic;
signal \N__27189\ : std_logic;
signal \N__27180\ : std_logic;
signal \N__27169\ : std_logic;
signal \N__27166\ : std_logic;
signal \N__27163\ : std_logic;
signal \N__27162\ : std_logic;
signal \N__27161\ : std_logic;
signal \N__27160\ : std_logic;
signal \N__27159\ : std_logic;
signal \N__27156\ : std_logic;
signal \N__27153\ : std_logic;
signal \N__27148\ : std_logic;
signal \N__27145\ : std_logic;
signal \N__27142\ : std_logic;
signal \N__27139\ : std_logic;
signal \N__27130\ : std_logic;
signal \N__27127\ : std_logic;
signal \N__27126\ : std_logic;
signal \N__27123\ : std_logic;
signal \N__27120\ : std_logic;
signal \N__27119\ : std_logic;
signal \N__27118\ : std_logic;
signal \N__27115\ : std_logic;
signal \N__27112\ : std_logic;
signal \N__27109\ : std_logic;
signal \N__27106\ : std_logic;
signal \N__27103\ : std_logic;
signal \N__27100\ : std_logic;
signal \N__27091\ : std_logic;
signal \N__27090\ : std_logic;
signal \N__27089\ : std_logic;
signal \N__27086\ : std_logic;
signal \N__27085\ : std_logic;
signal \N__27082\ : std_logic;
signal \N__27081\ : std_logic;
signal \N__27078\ : std_logic;
signal \N__27075\ : std_logic;
signal \N__27068\ : std_logic;
signal \N__27065\ : std_logic;
signal \N__27062\ : std_logic;
signal \N__27059\ : std_logic;
signal \N__27052\ : std_logic;
signal \N__27051\ : std_logic;
signal \N__27050\ : std_logic;
signal \N__27047\ : std_logic;
signal \N__27046\ : std_logic;
signal \N__27045\ : std_logic;
signal \N__27044\ : std_logic;
signal \N__27043\ : std_logic;
signal \N__27040\ : std_logic;
signal \N__27037\ : std_logic;
signal \N__27034\ : std_logic;
signal \N__27025\ : std_logic;
signal \N__27016\ : std_logic;
signal \N__27013\ : std_logic;
signal \N__27010\ : std_logic;
signal \N__27007\ : std_logic;
signal \N__27006\ : std_logic;
signal \N__27003\ : std_logic;
signal \N__27002\ : std_logic;
signal \N__26995\ : std_logic;
signal \N__26992\ : std_logic;
signal \N__26989\ : std_logic;
signal \N__26988\ : std_logic;
signal \N__26983\ : std_logic;
signal \N__26980\ : std_logic;
signal \N__26977\ : std_logic;
signal \N__26974\ : std_logic;
signal \N__26971\ : std_logic;
signal \N__26970\ : std_logic;
signal \N__26969\ : std_logic;
signal \N__26962\ : std_logic;
signal \N__26961\ : std_logic;
signal \N__26960\ : std_logic;
signal \N__26957\ : std_logic;
signal \N__26954\ : std_logic;
signal \N__26951\ : std_logic;
signal \N__26950\ : std_logic;
signal \N__26947\ : std_logic;
signal \N__26944\ : std_logic;
signal \N__26939\ : std_logic;
signal \N__26932\ : std_logic;
signal \N__26929\ : std_logic;
signal \N__26926\ : std_logic;
signal \N__26923\ : std_logic;
signal \N__26920\ : std_logic;
signal \N__26919\ : std_logic;
signal \N__26918\ : std_logic;
signal \N__26915\ : std_logic;
signal \N__26910\ : std_logic;
signal \N__26907\ : std_logic;
signal \N__26902\ : std_logic;
signal \N__26899\ : std_logic;
signal \N__26896\ : std_logic;
signal \N__26893\ : std_logic;
signal \N__26890\ : std_logic;
signal \N__26887\ : std_logic;
signal \N__26886\ : std_logic;
signal \N__26883\ : std_logic;
signal \N__26880\ : std_logic;
signal \N__26877\ : std_logic;
signal \N__26874\ : std_logic;
signal \N__26873\ : std_logic;
signal \N__26872\ : std_logic;
signal \N__26871\ : std_logic;
signal \N__26870\ : std_logic;
signal \N__26867\ : std_logic;
signal \N__26864\ : std_logic;
signal \N__26861\ : std_logic;
signal \N__26854\ : std_logic;
signal \N__26851\ : std_logic;
signal \N__26846\ : std_logic;
signal \N__26839\ : std_logic;
signal \N__26836\ : std_logic;
signal \N__26833\ : std_logic;
signal \N__26832\ : std_logic;
signal \N__26831\ : std_logic;
signal \N__26828\ : std_logic;
signal \N__26825\ : std_logic;
signal \N__26824\ : std_logic;
signal \N__26821\ : std_logic;
signal \N__26818\ : std_logic;
signal \N__26815\ : std_logic;
signal \N__26810\ : std_logic;
signal \N__26807\ : std_logic;
signal \N__26800\ : std_logic;
signal \N__26797\ : std_logic;
signal \N__26796\ : std_logic;
signal \N__26795\ : std_logic;
signal \N__26794\ : std_logic;
signal \N__26791\ : std_logic;
signal \N__26786\ : std_logic;
signal \N__26785\ : std_logic;
signal \N__26784\ : std_logic;
signal \N__26781\ : std_logic;
signal \N__26778\ : std_logic;
signal \N__26775\ : std_logic;
signal \N__26770\ : std_logic;
signal \N__26761\ : std_logic;
signal \N__26760\ : std_logic;
signal \N__26757\ : std_logic;
signal \N__26754\ : std_logic;
signal \N__26749\ : std_logic;
signal \N__26748\ : std_logic;
signal \N__26745\ : std_logic;
signal \N__26742\ : std_logic;
signal \N__26739\ : std_logic;
signal \N__26734\ : std_logic;
signal \N__26733\ : std_logic;
signal \N__26732\ : std_logic;
signal \N__26731\ : std_logic;
signal \N__26730\ : std_logic;
signal \N__26729\ : std_logic;
signal \N__26726\ : std_logic;
signal \N__26719\ : std_logic;
signal \N__26714\ : std_logic;
signal \N__26713\ : std_logic;
signal \N__26710\ : std_logic;
signal \N__26705\ : std_logic;
signal \N__26702\ : std_logic;
signal \N__26699\ : std_logic;
signal \N__26696\ : std_logic;
signal \N__26693\ : std_logic;
signal \N__26688\ : std_logic;
signal \N__26685\ : std_logic;
signal \N__26680\ : std_logic;
signal \N__26679\ : std_logic;
signal \N__26678\ : std_logic;
signal \N__26677\ : std_logic;
signal \N__26676\ : std_logic;
signal \N__26675\ : std_logic;
signal \N__26668\ : std_logic;
signal \N__26667\ : std_logic;
signal \N__26662\ : std_logic;
signal \N__26659\ : std_logic;
signal \N__26656\ : std_logic;
signal \N__26653\ : std_logic;
signal \N__26646\ : std_logic;
signal \N__26641\ : std_logic;
signal \N__26638\ : std_logic;
signal \N__26637\ : std_logic;
signal \N__26636\ : std_logic;
signal \N__26631\ : std_logic;
signal \N__26628\ : std_logic;
signal \N__26623\ : std_logic;
signal \N__26622\ : std_logic;
signal \N__26621\ : std_logic;
signal \N__26620\ : std_logic;
signal \N__26611\ : std_logic;
signal \N__26608\ : std_logic;
signal \N__26605\ : std_logic;
signal \N__26602\ : std_logic;
signal \N__26599\ : std_logic;
signal \N__26596\ : std_logic;
signal \N__26593\ : std_logic;
signal \N__26590\ : std_logic;
signal \N__26587\ : std_logic;
signal \N__26584\ : std_logic;
signal \N__26583\ : std_logic;
signal \N__26580\ : std_logic;
signal \N__26577\ : std_logic;
signal \N__26572\ : std_logic;
signal \N__26569\ : std_logic;
signal \N__26566\ : std_logic;
signal \N__26565\ : std_logic;
signal \N__26562\ : std_logic;
signal \N__26559\ : std_logic;
signal \N__26554\ : std_logic;
signal \N__26551\ : std_logic;
signal \N__26548\ : std_logic;
signal \N__26545\ : std_logic;
signal \N__26542\ : std_logic;
signal \N__26541\ : std_logic;
signal \N__26540\ : std_logic;
signal \N__26537\ : std_logic;
signal \N__26532\ : std_logic;
signal \N__26527\ : std_logic;
signal \N__26526\ : std_logic;
signal \N__26523\ : std_logic;
signal \N__26520\ : std_logic;
signal \N__26515\ : std_logic;
signal \N__26512\ : std_logic;
signal \N__26511\ : std_logic;
signal \N__26510\ : std_logic;
signal \N__26509\ : std_logic;
signal \N__26504\ : std_logic;
signal \N__26503\ : std_logic;
signal \N__26502\ : std_logic;
signal \N__26501\ : std_logic;
signal \N__26500\ : std_logic;
signal \N__26497\ : std_logic;
signal \N__26496\ : std_logic;
signal \N__26495\ : std_logic;
signal \N__26492\ : std_logic;
signal \N__26491\ : std_logic;
signal \N__26490\ : std_logic;
signal \N__26487\ : std_logic;
signal \N__26486\ : std_logic;
signal \N__26483\ : std_logic;
signal \N__26478\ : std_logic;
signal \N__26469\ : std_logic;
signal \N__26466\ : std_logic;
signal \N__26461\ : std_logic;
signal \N__26458\ : std_logic;
signal \N__26455\ : std_logic;
signal \N__26440\ : std_logic;
signal \N__26439\ : std_logic;
signal \N__26434\ : std_logic;
signal \N__26431\ : std_logic;
signal \N__26428\ : std_logic;
signal \N__26427\ : std_logic;
signal \N__26426\ : std_logic;
signal \N__26425\ : std_logic;
signal \N__26418\ : std_logic;
signal \N__26417\ : std_logic;
signal \N__26414\ : std_logic;
signal \N__26411\ : std_logic;
signal \N__26410\ : std_logic;
signal \N__26409\ : std_logic;
signal \N__26408\ : std_logic;
signal \N__26407\ : std_logic;
signal \N__26406\ : std_logic;
signal \N__26403\ : std_logic;
signal \N__26402\ : std_logic;
signal \N__26401\ : std_logic;
signal \N__26398\ : std_logic;
signal \N__26395\ : std_logic;
signal \N__26386\ : std_logic;
signal \N__26383\ : std_logic;
signal \N__26376\ : std_logic;
signal \N__26365\ : std_logic;
signal \N__26362\ : std_logic;
signal \N__26359\ : std_logic;
signal \N__26356\ : std_logic;
signal \N__26355\ : std_logic;
signal \N__26354\ : std_logic;
signal \N__26351\ : std_logic;
signal \N__26346\ : std_logic;
signal \N__26341\ : std_logic;
signal \N__26338\ : std_logic;
signal \N__26337\ : std_logic;
signal \N__26336\ : std_logic;
signal \N__26335\ : std_logic;
signal \N__26334\ : std_logic;
signal \N__26333\ : std_logic;
signal \N__26332\ : std_logic;
signal \N__26331\ : std_logic;
signal \N__26328\ : std_logic;
signal \N__26321\ : std_logic;
signal \N__26318\ : std_logic;
signal \N__26317\ : std_logic;
signal \N__26310\ : std_logic;
signal \N__26305\ : std_logic;
signal \N__26302\ : std_logic;
signal \N__26301\ : std_logic;
signal \N__26300\ : std_logic;
signal \N__26299\ : std_logic;
signal \N__26298\ : std_logic;
signal \N__26297\ : std_logic;
signal \N__26294\ : std_logic;
signal \N__26293\ : std_logic;
signal \N__26292\ : std_logic;
signal \N__26289\ : std_logic;
signal \N__26284\ : std_logic;
signal \N__26273\ : std_logic;
signal \N__26266\ : std_logic;
signal \N__26257\ : std_logic;
signal \N__26254\ : std_logic;
signal \N__26251\ : std_logic;
signal \N__26248\ : std_logic;
signal \N__26245\ : std_logic;
signal \N__26242\ : std_logic;
signal \N__26239\ : std_logic;
signal \N__26236\ : std_logic;
signal \N__26233\ : std_logic;
signal \N__26230\ : std_logic;
signal \N__26229\ : std_logic;
signal \N__26226\ : std_logic;
signal \N__26225\ : std_logic;
signal \N__26224\ : std_logic;
signal \N__26223\ : std_logic;
signal \N__26220\ : std_logic;
signal \N__26217\ : std_logic;
signal \N__26214\ : std_logic;
signal \N__26209\ : std_logic;
signal \N__26206\ : std_logic;
signal \N__26197\ : std_logic;
signal \N__26194\ : std_logic;
signal \N__26193\ : std_logic;
signal \N__26192\ : std_logic;
signal \N__26189\ : std_logic;
signal \N__26188\ : std_logic;
signal \N__26185\ : std_logic;
signal \N__26182\ : std_logic;
signal \N__26179\ : std_logic;
signal \N__26176\ : std_logic;
signal \N__26171\ : std_logic;
signal \N__26166\ : std_logic;
signal \N__26161\ : std_logic;
signal \N__26158\ : std_logic;
signal \N__26157\ : std_logic;
signal \N__26156\ : std_logic;
signal \N__26153\ : std_logic;
signal \N__26152\ : std_logic;
signal \N__26151\ : std_logic;
signal \N__26150\ : std_logic;
signal \N__26149\ : std_logic;
signal \N__26148\ : std_logic;
signal \N__26147\ : std_logic;
signal \N__26146\ : std_logic;
signal \N__26145\ : std_logic;
signal \N__26144\ : std_logic;
signal \N__26143\ : std_logic;
signal \N__26138\ : std_logic;
signal \N__26135\ : std_logic;
signal \N__26130\ : std_logic;
signal \N__26127\ : std_logic;
signal \N__26124\ : std_logic;
signal \N__26121\ : std_logic;
signal \N__26118\ : std_logic;
signal \N__26115\ : std_logic;
signal \N__26110\ : std_logic;
signal \N__26107\ : std_logic;
signal \N__26106\ : std_logic;
signal \N__26105\ : std_logic;
signal \N__26104\ : std_logic;
signal \N__26103\ : std_logic;
signal \N__26102\ : std_logic;
signal \N__26101\ : std_logic;
signal \N__26100\ : std_logic;
signal \N__26099\ : std_logic;
signal \N__26098\ : std_logic;
signal \N__26097\ : std_logic;
signal \N__26096\ : std_logic;
signal \N__26095\ : std_logic;
signal \N__26094\ : std_logic;
signal \N__26093\ : std_logic;
signal \N__26092\ : std_logic;
signal \N__26091\ : std_logic;
signal \N__26090\ : std_logic;
signal \N__26089\ : std_logic;
signal \N__26088\ : std_logic;
signal \N__26087\ : std_logic;
signal \N__26086\ : std_logic;
signal \N__26085\ : std_logic;
signal \N__26084\ : std_logic;
signal \N__26083\ : std_logic;
signal \N__26082\ : std_logic;
signal \N__26081\ : std_logic;
signal \N__26080\ : std_logic;
signal \N__26079\ : std_logic;
signal \N__26078\ : std_logic;
signal \N__26077\ : std_logic;
signal \N__26076\ : std_logic;
signal \N__26075\ : std_logic;
signal \N__26074\ : std_logic;
signal \N__26073\ : std_logic;
signal \N__26072\ : std_logic;
signal \N__26071\ : std_logic;
signal \N__26070\ : std_logic;
signal \N__26069\ : std_logic;
signal \N__26068\ : std_logic;
signal \N__26067\ : std_logic;
signal \N__26066\ : std_logic;
signal \N__26065\ : std_logic;
signal \N__26064\ : std_logic;
signal \N__26063\ : std_logic;
signal \N__26060\ : std_logic;
signal \N__26057\ : std_logic;
signal \N__26054\ : std_logic;
signal \N__26051\ : std_logic;
signal \N__26050\ : std_logic;
signal \N__26049\ : std_logic;
signal \N__26048\ : std_logic;
signal \N__26047\ : std_logic;
signal \N__26046\ : std_logic;
signal \N__26045\ : std_logic;
signal \N__26044\ : std_logic;
signal \N__26043\ : std_logic;
signal \N__26042\ : std_logic;
signal \N__26041\ : std_logic;
signal \N__26040\ : std_logic;
signal \N__26039\ : std_logic;
signal \N__26038\ : std_logic;
signal \N__26037\ : std_logic;
signal \N__26034\ : std_logic;
signal \N__26031\ : std_logic;
signal \N__26028\ : std_logic;
signal \N__26025\ : std_logic;
signal \N__26022\ : std_logic;
signal \N__26019\ : std_logic;
signal \N__25882\ : std_logic;
signal \N__25879\ : std_logic;
signal \N__25876\ : std_logic;
signal \N__25875\ : std_logic;
signal \N__25870\ : std_logic;
signal \N__25867\ : std_logic;
signal \N__25866\ : std_logic;
signal \N__25865\ : std_logic;
signal \N__25862\ : std_logic;
signal \N__25857\ : std_logic;
signal \N__25852\ : std_logic;
signal \N__25851\ : std_logic;
signal \N__25848\ : std_logic;
signal \N__25845\ : std_logic;
signal \N__25844\ : std_logic;
signal \N__25843\ : std_logic;
signal \N__25840\ : std_logic;
signal \N__25837\ : std_logic;
signal \N__25834\ : std_logic;
signal \N__25831\ : std_logic;
signal \N__25828\ : std_logic;
signal \N__25823\ : std_logic;
signal \N__25816\ : std_logic;
signal \N__25813\ : std_logic;
signal \N__25810\ : std_logic;
signal \N__25809\ : std_logic;
signal \N__25806\ : std_logic;
signal \N__25803\ : std_logic;
signal \N__25802\ : std_logic;
signal \N__25799\ : std_logic;
signal \N__25796\ : std_logic;
signal \N__25793\ : std_logic;
signal \N__25788\ : std_logic;
signal \N__25783\ : std_logic;
signal \N__25780\ : std_logic;
signal \N__25779\ : std_logic;
signal \N__25776\ : std_logic;
signal \N__25775\ : std_logic;
signal \N__25772\ : std_logic;
signal \N__25769\ : std_logic;
signal \N__25766\ : std_logic;
signal \N__25763\ : std_logic;
signal \N__25760\ : std_logic;
signal \N__25753\ : std_logic;
signal \N__25750\ : std_logic;
signal \N__25747\ : std_logic;
signal \N__25744\ : std_logic;
signal \N__25741\ : std_logic;
signal \N__25738\ : std_logic;
signal \N__25735\ : std_logic;
signal \N__25732\ : std_logic;
signal \N__25729\ : std_logic;
signal \N__25728\ : std_logic;
signal \N__25725\ : std_logic;
signal \N__25724\ : std_logic;
signal \N__25721\ : std_logic;
signal \N__25718\ : std_logic;
signal \N__25715\ : std_logic;
signal \N__25708\ : std_logic;
signal \N__25705\ : std_logic;
signal \N__25702\ : std_logic;
signal \N__25699\ : std_logic;
signal \N__25696\ : std_logic;
signal \N__25693\ : std_logic;
signal \N__25690\ : std_logic;
signal \N__25687\ : std_logic;
signal \N__25684\ : std_logic;
signal \N__25683\ : std_logic;
signal \N__25682\ : std_logic;
signal \N__25677\ : std_logic;
signal \N__25674\ : std_logic;
signal \N__25671\ : std_logic;
signal \N__25668\ : std_logic;
signal \N__25665\ : std_logic;
signal \N__25660\ : std_logic;
signal \N__25659\ : std_logic;
signal \N__25654\ : std_logic;
signal \N__25651\ : std_logic;
signal \N__25648\ : std_logic;
signal \N__25645\ : std_logic;
signal \N__25642\ : std_logic;
signal \N__25639\ : std_logic;
signal \N__25636\ : std_logic;
signal \N__25633\ : std_logic;
signal \N__25630\ : std_logic;
signal \N__25629\ : std_logic;
signal \N__25626\ : std_logic;
signal \N__25625\ : std_logic;
signal \N__25622\ : std_logic;
signal \N__25619\ : std_logic;
signal \N__25616\ : std_logic;
signal \N__25609\ : std_logic;
signal \N__25606\ : std_logic;
signal \N__25603\ : std_logic;
signal \N__25600\ : std_logic;
signal \N__25597\ : std_logic;
signal \N__25594\ : std_logic;
signal \N__25591\ : std_logic;
signal \N__25590\ : std_logic;
signal \N__25587\ : std_logic;
signal \N__25586\ : std_logic;
signal \N__25583\ : std_logic;
signal \N__25580\ : std_logic;
signal \N__25577\ : std_logic;
signal \N__25570\ : std_logic;
signal \N__25567\ : std_logic;
signal \N__25566\ : std_logic;
signal \N__25565\ : std_logic;
signal \N__25558\ : std_logic;
signal \N__25555\ : std_logic;
signal \N__25552\ : std_logic;
signal \N__25551\ : std_logic;
signal \N__25546\ : std_logic;
signal \N__25543\ : std_logic;
signal \N__25540\ : std_logic;
signal \N__25537\ : std_logic;
signal \N__25534\ : std_logic;
signal \N__25533\ : std_logic;
signal \N__25530\ : std_logic;
signal \N__25527\ : std_logic;
signal \N__25526\ : std_logic;
signal \N__25523\ : std_logic;
signal \N__25520\ : std_logic;
signal \N__25517\ : std_logic;
signal \N__25514\ : std_logic;
signal \N__25511\ : std_logic;
signal \N__25504\ : std_logic;
signal \N__25501\ : std_logic;
signal \N__25498\ : std_logic;
signal \N__25495\ : std_logic;
signal \N__25492\ : std_logic;
signal \N__25491\ : std_logic;
signal \N__25490\ : std_logic;
signal \N__25489\ : std_logic;
signal \N__25486\ : std_logic;
signal \N__25479\ : std_logic;
signal \N__25478\ : std_logic;
signal \N__25477\ : std_logic;
signal \N__25474\ : std_logic;
signal \N__25471\ : std_logic;
signal \N__25466\ : std_logic;
signal \N__25461\ : std_logic;
signal \N__25456\ : std_logic;
signal \N__25453\ : std_logic;
signal \N__25452\ : std_logic;
signal \N__25447\ : std_logic;
signal \N__25444\ : std_logic;
signal \N__25441\ : std_logic;
signal \N__25438\ : std_logic;
signal \N__25435\ : std_logic;
signal \N__25432\ : std_logic;
signal \N__25429\ : std_logic;
signal \N__25428\ : std_logic;
signal \N__25427\ : std_logic;
signal \N__25426\ : std_logic;
signal \N__25425\ : std_logic;
signal \N__25424\ : std_logic;
signal \N__25423\ : std_logic;
signal \N__25408\ : std_logic;
signal \N__25405\ : std_logic;
signal \N__25402\ : std_logic;
signal \N__25399\ : std_logic;
signal \N__25398\ : std_logic;
signal \N__25397\ : std_logic;
signal \N__25396\ : std_logic;
signal \N__25395\ : std_logic;
signal \N__25394\ : std_logic;
signal \N__25391\ : std_logic;
signal \N__25386\ : std_logic;
signal \N__25381\ : std_logic;
signal \N__25378\ : std_logic;
signal \N__25377\ : std_logic;
signal \N__25376\ : std_logic;
signal \N__25375\ : std_logic;
signal \N__25374\ : std_logic;
signal \N__25373\ : std_logic;
signal \N__25372\ : std_logic;
signal \N__25363\ : std_logic;
signal \N__25360\ : std_logic;
signal \N__25357\ : std_logic;
signal \N__25350\ : std_logic;
signal \N__25347\ : std_logic;
signal \N__25346\ : std_logic;
signal \N__25345\ : std_logic;
signal \N__25344\ : std_logic;
signal \N__25341\ : std_logic;
signal \N__25334\ : std_logic;
signal \N__25331\ : std_logic;
signal \N__25324\ : std_logic;
signal \N__25315\ : std_logic;
signal \N__25314\ : std_logic;
signal \N__25313\ : std_logic;
signal \N__25308\ : std_logic;
signal \N__25305\ : std_logic;
signal \N__25304\ : std_logic;
signal \N__25303\ : std_logic;
signal \N__25302\ : std_logic;
signal \N__25301\ : std_logic;
signal \N__25300\ : std_logic;
signal \N__25297\ : std_logic;
signal \N__25294\ : std_logic;
signal \N__25291\ : std_logic;
signal \N__25288\ : std_logic;
signal \N__25283\ : std_logic;
signal \N__25280\ : std_logic;
signal \N__25279\ : std_logic;
signal \N__25274\ : std_logic;
signal \N__25273\ : std_logic;
signal \N__25272\ : std_logic;
signal \N__25269\ : std_logic;
signal \N__25266\ : std_logic;
signal \N__25261\ : std_logic;
signal \N__25260\ : std_logic;
signal \N__25257\ : std_logic;
signal \N__25254\ : std_logic;
signal \N__25251\ : std_logic;
signal \N__25248\ : std_logic;
signal \N__25241\ : std_logic;
signal \N__25238\ : std_logic;
signal \N__25225\ : std_logic;
signal \N__25222\ : std_logic;
signal \N__25219\ : std_logic;
signal \N__25216\ : std_logic;
signal \N__25213\ : std_logic;
signal \N__25212\ : std_logic;
signal \N__25211\ : std_logic;
signal \N__25210\ : std_logic;
signal \N__25201\ : std_logic;
signal \N__25200\ : std_logic;
signal \N__25199\ : std_logic;
signal \N__25196\ : std_logic;
signal \N__25193\ : std_logic;
signal \N__25190\ : std_logic;
signal \N__25185\ : std_logic;
signal \N__25180\ : std_logic;
signal \N__25179\ : std_logic;
signal \N__25176\ : std_logic;
signal \N__25173\ : std_logic;
signal \N__25170\ : std_logic;
signal \N__25167\ : std_logic;
signal \N__25162\ : std_logic;
signal \N__25161\ : std_logic;
signal \N__25160\ : std_logic;
signal \N__25157\ : std_logic;
signal \N__25152\ : std_logic;
signal \N__25147\ : std_logic;
signal \N__25146\ : std_logic;
signal \N__25143\ : std_logic;
signal \N__25140\ : std_logic;
signal \N__25137\ : std_logic;
signal \N__25134\ : std_logic;
signal \N__25133\ : std_logic;
signal \N__25132\ : std_logic;
signal \N__25131\ : std_logic;
signal \N__25126\ : std_logic;
signal \N__25119\ : std_logic;
signal \N__25114\ : std_logic;
signal \N__25111\ : std_logic;
signal \N__25110\ : std_logic;
signal \N__25109\ : std_logic;
signal \N__25108\ : std_logic;
signal \N__25105\ : std_logic;
signal \N__25100\ : std_logic;
signal \N__25097\ : std_logic;
signal \N__25092\ : std_logic;
signal \N__25089\ : std_logic;
signal \N__25088\ : std_logic;
signal \N__25085\ : std_logic;
signal \N__25082\ : std_logic;
signal \N__25079\ : std_logic;
signal \N__25076\ : std_logic;
signal \N__25069\ : std_logic;
signal \N__25066\ : std_logic;
signal \N__25063\ : std_logic;
signal \N__25062\ : std_logic;
signal \N__25061\ : std_logic;
signal \N__25058\ : std_logic;
signal \N__25053\ : std_logic;
signal \N__25048\ : std_logic;
signal \N__25047\ : std_logic;
signal \N__25046\ : std_logic;
signal \N__25045\ : std_logic;
signal \N__25042\ : std_logic;
signal \N__25041\ : std_logic;
signal \N__25040\ : std_logic;
signal \N__25039\ : std_logic;
signal \N__25036\ : std_logic;
signal \N__25033\ : std_logic;
signal \N__25026\ : std_logic;
signal \N__25025\ : std_logic;
signal \N__25024\ : std_logic;
signal \N__25023\ : std_logic;
signal \N__25022\ : std_logic;
signal \N__25021\ : std_logic;
signal \N__25020\ : std_logic;
signal \N__25019\ : std_logic;
signal \N__25016\ : std_logic;
signal \N__25013\ : std_logic;
signal \N__25012\ : std_logic;
signal \N__25011\ : std_logic;
signal \N__25010\ : std_logic;
signal \N__25009\ : std_logic;
signal \N__25008\ : std_logic;
signal \N__25005\ : std_logic;
signal \N__25002\ : std_logic;
signal \N__24999\ : std_logic;
signal \N__24996\ : std_logic;
signal \N__24987\ : std_logic;
signal \N__24982\ : std_logic;
signal \N__24979\ : std_logic;
signal \N__24976\ : std_logic;
signal \N__24973\ : std_logic;
signal \N__24968\ : std_logic;
signal \N__24965\ : std_logic;
signal \N__24964\ : std_logic;
signal \N__24961\ : std_logic;
signal \N__24958\ : std_logic;
signal \N__24953\ : std_logic;
signal \N__24950\ : std_logic;
signal \N__24947\ : std_logic;
signal \N__24944\ : std_logic;
signal \N__24935\ : std_logic;
signal \N__24930\ : std_logic;
signal \N__24927\ : std_logic;
signal \N__24922\ : std_logic;
signal \N__24919\ : std_logic;
signal \N__24910\ : std_logic;
signal \N__24901\ : std_logic;
signal \N__24900\ : std_logic;
signal \N__24899\ : std_logic;
signal \N__24898\ : std_logic;
signal \N__24897\ : std_logic;
signal \N__24894\ : std_logic;
signal \N__24891\ : std_logic;
signal \N__24890\ : std_logic;
signal \N__24889\ : std_logic;
signal \N__24888\ : std_logic;
signal \N__24887\ : std_logic;
signal \N__24886\ : std_logic;
signal \N__24885\ : std_logic;
signal \N__24882\ : std_logic;
signal \N__24879\ : std_logic;
signal \N__24878\ : std_logic;
signal \N__24875\ : std_logic;
signal \N__24874\ : std_logic;
signal \N__24871\ : std_logic;
signal \N__24868\ : std_logic;
signal \N__24865\ : std_logic;
signal \N__24864\ : std_logic;
signal \N__24863\ : std_logic;
signal \N__24862\ : std_logic;
signal \N__24861\ : std_logic;
signal \N__24856\ : std_logic;
signal \N__24849\ : std_logic;
signal \N__24844\ : std_logic;
signal \N__24841\ : std_logic;
signal \N__24838\ : std_logic;
signal \N__24835\ : std_logic;
signal \N__24830\ : std_logic;
signal \N__24827\ : std_logic;
signal \N__24824\ : std_logic;
signal \N__24819\ : std_logic;
signal \N__24816\ : std_logic;
signal \N__24815\ : std_logic;
signal \N__24814\ : std_logic;
signal \N__24813\ : std_logic;
signal \N__24810\ : std_logic;
signal \N__24807\ : std_logic;
signal \N__24804\ : std_logic;
signal \N__24803\ : std_logic;
signal \N__24802\ : std_logic;
signal \N__24797\ : std_logic;
signal \N__24790\ : std_logic;
signal \N__24787\ : std_logic;
signal \N__24784\ : std_logic;
signal \N__24779\ : std_logic;
signal \N__24774\ : std_logic;
signal \N__24767\ : std_logic;
signal \N__24762\ : std_logic;
signal \N__24757\ : std_logic;
signal \N__24742\ : std_logic;
signal \N__24739\ : std_logic;
signal \N__24736\ : std_logic;
signal \N__24733\ : std_logic;
signal \N__24730\ : std_logic;
signal \N__24727\ : std_logic;
signal \N__24726\ : std_logic;
signal \N__24725\ : std_logic;
signal \N__24720\ : std_logic;
signal \N__24717\ : std_logic;
signal \N__24714\ : std_logic;
signal \N__24711\ : std_logic;
signal \N__24706\ : std_logic;
signal \N__24705\ : std_logic;
signal \N__24704\ : std_logic;
signal \N__24703\ : std_logic;
signal \N__24702\ : std_logic;
signal \N__24699\ : std_logic;
signal \N__24696\ : std_logic;
signal \N__24695\ : std_logic;
signal \N__24690\ : std_logic;
signal \N__24689\ : std_logic;
signal \N__24688\ : std_logic;
signal \N__24687\ : std_logic;
signal \N__24686\ : std_logic;
signal \N__24685\ : std_logic;
signal \N__24684\ : std_logic;
signal \N__24683\ : std_logic;
signal \N__24682\ : std_logic;
signal \N__24681\ : std_logic;
signal \N__24680\ : std_logic;
signal \N__24679\ : std_logic;
signal \N__24678\ : std_logic;
signal \N__24677\ : std_logic;
signal \N__24676\ : std_logic;
signal \N__24675\ : std_logic;
signal \N__24674\ : std_logic;
signal \N__24673\ : std_logic;
signal \N__24672\ : std_logic;
signal \N__24671\ : std_logic;
signal \N__24670\ : std_logic;
signal \N__24669\ : std_logic;
signal \N__24666\ : std_logic;
signal \N__24663\ : std_logic;
signal \N__24660\ : std_logic;
signal \N__24657\ : std_logic;
signal \N__24654\ : std_logic;
signal \N__24651\ : std_logic;
signal \N__24644\ : std_logic;
signal \N__24637\ : std_logic;
signal \N__24634\ : std_logic;
signal \N__24631\ : std_logic;
signal \N__24628\ : std_logic;
signal \N__24627\ : std_logic;
signal \N__24626\ : std_logic;
signal \N__24623\ : std_logic;
signal \N__24618\ : std_logic;
signal \N__24615\ : std_logic;
signal \N__24606\ : std_logic;
signal \N__24599\ : std_logic;
signal \N__24596\ : std_logic;
signal \N__24591\ : std_logic;
signal \N__24584\ : std_logic;
signal \N__24579\ : std_logic;
signal \N__24578\ : std_logic;
signal \N__24577\ : std_logic;
signal \N__24574\ : std_logic;
signal \N__24569\ : std_logic;
signal \N__24564\ : std_logic;
signal \N__24557\ : std_logic;
signal \N__24550\ : std_logic;
signal \N__24547\ : std_logic;
signal \N__24542\ : std_logic;
signal \N__24537\ : std_logic;
signal \N__24532\ : std_logic;
signal \N__24525\ : std_logic;
signal \N__24514\ : std_logic;
signal \N__24513\ : std_logic;
signal \N__24512\ : std_logic;
signal \N__24509\ : std_logic;
signal \N__24504\ : std_logic;
signal \N__24499\ : std_logic;
signal \N__24496\ : std_logic;
signal \N__24495\ : std_logic;
signal \N__24490\ : std_logic;
signal \N__24487\ : std_logic;
signal \N__24484\ : std_logic;
signal \N__24481\ : std_logic;
signal \N__24478\ : std_logic;
signal \N__24477\ : std_logic;
signal \N__24476\ : std_logic;
signal \N__24475\ : std_logic;
signal \N__24472\ : std_logic;
signal \N__24469\ : std_logic;
signal \N__24466\ : std_logic;
signal \N__24463\ : std_logic;
signal \N__24460\ : std_logic;
signal \N__24457\ : std_logic;
signal \N__24448\ : std_logic;
signal \N__24447\ : std_logic;
signal \N__24446\ : std_logic;
signal \N__24445\ : std_logic;
signal \N__24444\ : std_logic;
signal \N__24443\ : std_logic;
signal \N__24442\ : std_logic;
signal \N__24441\ : std_logic;
signal \N__24440\ : std_logic;
signal \N__24437\ : std_logic;
signal \N__24434\ : std_logic;
signal \N__24429\ : std_logic;
signal \N__24426\ : std_logic;
signal \N__24423\ : std_logic;
signal \N__24418\ : std_logic;
signal \N__24417\ : std_logic;
signal \N__24416\ : std_logic;
signal \N__24415\ : std_logic;
signal \N__24414\ : std_logic;
signal \N__24411\ : std_logic;
signal \N__24408\ : std_logic;
signal \N__24401\ : std_logic;
signal \N__24398\ : std_logic;
signal \N__24395\ : std_logic;
signal \N__24392\ : std_logic;
signal \N__24387\ : std_logic;
signal \N__24384\ : std_logic;
signal \N__24379\ : std_logic;
signal \N__24376\ : std_logic;
signal \N__24371\ : std_logic;
signal \N__24358\ : std_logic;
signal \N__24357\ : std_logic;
signal \N__24356\ : std_logic;
signal \N__24351\ : std_logic;
signal \N__24348\ : std_logic;
signal \N__24347\ : std_logic;
signal \N__24344\ : std_logic;
signal \N__24341\ : std_logic;
signal \N__24340\ : std_logic;
signal \N__24337\ : std_logic;
signal \N__24332\ : std_logic;
signal \N__24329\ : std_logic;
signal \N__24322\ : std_logic;
signal \N__24321\ : std_logic;
signal \N__24320\ : std_logic;
signal \N__24317\ : std_logic;
signal \N__24314\ : std_logic;
signal \N__24311\ : std_logic;
signal \N__24310\ : std_logic;
signal \N__24309\ : std_logic;
signal \N__24308\ : std_logic;
signal \N__24301\ : std_logic;
signal \N__24300\ : std_logic;
signal \N__24297\ : std_logic;
signal \N__24296\ : std_logic;
signal \N__24295\ : std_logic;
signal \N__24294\ : std_logic;
signal \N__24291\ : std_logic;
signal \N__24288\ : std_logic;
signal \N__24285\ : std_logic;
signal \N__24282\ : std_logic;
signal \N__24275\ : std_logic;
signal \N__24272\ : std_logic;
signal \N__24271\ : std_logic;
signal \N__24270\ : std_logic;
signal \N__24267\ : std_logic;
signal \N__24266\ : std_logic;
signal \N__24263\ : std_logic;
signal \N__24260\ : std_logic;
signal \N__24255\ : std_logic;
signal \N__24252\ : std_logic;
signal \N__24247\ : std_logic;
signal \N__24244\ : std_logic;
signal \N__24241\ : std_logic;
signal \N__24238\ : std_logic;
signal \N__24235\ : std_logic;
signal \N__24230\ : std_logic;
signal \N__24217\ : std_logic;
signal \N__24214\ : std_logic;
signal \N__24211\ : std_logic;
signal \N__24208\ : std_logic;
signal \N__24207\ : std_logic;
signal \N__24206\ : std_logic;
signal \N__24203\ : std_logic;
signal \N__24200\ : std_logic;
signal \N__24197\ : std_logic;
signal \N__24194\ : std_logic;
signal \N__24191\ : std_logic;
signal \N__24188\ : std_logic;
signal \N__24185\ : std_logic;
signal \N__24178\ : std_logic;
signal \N__24177\ : std_logic;
signal \N__24176\ : std_logic;
signal \N__24173\ : std_logic;
signal \N__24172\ : std_logic;
signal \N__24169\ : std_logic;
signal \N__24168\ : std_logic;
signal \N__24165\ : std_logic;
signal \N__24162\ : std_logic;
signal \N__24159\ : std_logic;
signal \N__24158\ : std_logic;
signal \N__24157\ : std_logic;
signal \N__24150\ : std_logic;
signal \N__24145\ : std_logic;
signal \N__24140\ : std_logic;
signal \N__24133\ : std_logic;
signal \N__24130\ : std_logic;
signal \N__24127\ : std_logic;
signal \N__24126\ : std_logic;
signal \N__24123\ : std_logic;
signal \N__24122\ : std_logic;
signal \N__24121\ : std_logic;
signal \N__24120\ : std_logic;
signal \N__24113\ : std_logic;
signal \N__24110\ : std_logic;
signal \N__24107\ : std_logic;
signal \N__24104\ : std_logic;
signal \N__24101\ : std_logic;
signal \N__24098\ : std_logic;
signal \N__24095\ : std_logic;
signal \N__24088\ : std_logic;
signal \N__24085\ : std_logic;
signal \N__24084\ : std_logic;
signal \N__24081\ : std_logic;
signal \N__24078\ : std_logic;
signal \N__24073\ : std_logic;
signal \N__24072\ : std_logic;
signal \N__24069\ : std_logic;
signal \N__24068\ : std_logic;
signal \N__24061\ : std_logic;
signal \N__24058\ : std_logic;
signal \N__24057\ : std_logic;
signal \N__24056\ : std_logic;
signal \N__24055\ : std_logic;
signal \N__24054\ : std_logic;
signal \N__24053\ : std_logic;
signal \N__24052\ : std_logic;
signal \N__24047\ : std_logic;
signal \N__24044\ : std_logic;
signal \N__24035\ : std_logic;
signal \N__24028\ : std_logic;
signal \N__24025\ : std_logic;
signal \N__24022\ : std_logic;
signal \N__24019\ : std_logic;
signal \N__24016\ : std_logic;
signal \N__24013\ : std_logic;
signal \N__24012\ : std_logic;
signal \N__24011\ : std_logic;
signal \N__24008\ : std_logic;
signal \N__24007\ : std_logic;
signal \N__24006\ : std_logic;
signal \N__24005\ : std_logic;
signal \N__24004\ : std_logic;
signal \N__24003\ : std_logic;
signal \N__24000\ : std_logic;
signal \N__23997\ : std_logic;
signal \N__23994\ : std_logic;
signal \N__23991\ : std_logic;
signal \N__23988\ : std_logic;
signal \N__23985\ : std_logic;
signal \N__23982\ : std_logic;
signal \N__23977\ : std_logic;
signal \N__23976\ : std_logic;
signal \N__23973\ : std_logic;
signal \N__23972\ : std_logic;
signal \N__23969\ : std_logic;
signal \N__23966\ : std_logic;
signal \N__23963\ : std_logic;
signal \N__23960\ : std_logic;
signal \N__23955\ : std_logic;
signal \N__23952\ : std_logic;
signal \N__23949\ : std_logic;
signal \N__23946\ : std_logic;
signal \N__23937\ : std_logic;
signal \N__23934\ : std_logic;
signal \N__23923\ : std_logic;
signal \N__23920\ : std_logic;
signal \N__23917\ : std_logic;
signal \N__23914\ : std_logic;
signal \N__23913\ : std_logic;
signal \N__23910\ : std_logic;
signal \N__23907\ : std_logic;
signal \N__23902\ : std_logic;
signal \N__23899\ : std_logic;
signal \N__23898\ : std_logic;
signal \N__23895\ : std_logic;
signal \N__23892\ : std_logic;
signal \N__23889\ : std_logic;
signal \N__23886\ : std_logic;
signal \N__23883\ : std_logic;
signal \N__23880\ : std_logic;
signal \N__23877\ : std_logic;
signal \N__23874\ : std_logic;
signal \N__23869\ : std_logic;
signal \N__23866\ : std_logic;
signal \N__23863\ : std_logic;
signal \N__23860\ : std_logic;
signal \N__23857\ : std_logic;
signal \N__23856\ : std_logic;
signal \N__23855\ : std_logic;
signal \N__23854\ : std_logic;
signal \N__23851\ : std_logic;
signal \N__23846\ : std_logic;
signal \N__23843\ : std_logic;
signal \N__23836\ : std_logic;
signal \N__23833\ : std_logic;
signal \N__23832\ : std_logic;
signal \N__23831\ : std_logic;
signal \N__23828\ : std_logic;
signal \N__23827\ : std_logic;
signal \N__23826\ : std_logic;
signal \N__23825\ : std_logic;
signal \N__23824\ : std_logic;
signal \N__23819\ : std_logic;
signal \N__23818\ : std_logic;
signal \N__23817\ : std_logic;
signal \N__23816\ : std_logic;
signal \N__23815\ : std_logic;
signal \N__23814\ : std_logic;
signal \N__23813\ : std_logic;
signal \N__23812\ : std_logic;
signal \N__23807\ : std_logic;
signal \N__23804\ : std_logic;
signal \N__23799\ : std_logic;
signal \N__23798\ : std_logic;
signal \N__23795\ : std_logic;
signal \N__23792\ : std_logic;
signal \N__23789\ : std_logic;
signal \N__23786\ : std_logic;
signal \N__23785\ : std_logic;
signal \N__23784\ : std_logic;
signal \N__23781\ : std_logic;
signal \N__23778\ : std_logic;
signal \N__23777\ : std_logic;
signal \N__23776\ : std_logic;
signal \N__23775\ : std_logic;
signal \N__23772\ : std_logic;
signal \N__23769\ : std_logic;
signal \N__23764\ : std_logic;
signal \N__23761\ : std_logic;
signal \N__23758\ : std_logic;
signal \N__23749\ : std_logic;
signal \N__23744\ : std_logic;
signal \N__23741\ : std_logic;
signal \N__23738\ : std_logic;
signal \N__23731\ : std_logic;
signal \N__23724\ : std_logic;
signal \N__23721\ : std_logic;
signal \N__23716\ : std_logic;
signal \N__23709\ : std_logic;
signal \N__23704\ : std_logic;
signal \N__23699\ : std_logic;
signal \N__23696\ : std_logic;
signal \N__23693\ : std_logic;
signal \N__23686\ : std_logic;
signal \N__23685\ : std_logic;
signal \N__23682\ : std_logic;
signal \N__23679\ : std_logic;
signal \N__23674\ : std_logic;
signal \N__23671\ : std_logic;
signal \N__23670\ : std_logic;
signal \N__23665\ : std_logic;
signal \N__23662\ : std_logic;
signal \N__23659\ : std_logic;
signal \N__23656\ : std_logic;
signal \N__23655\ : std_logic;
signal \N__23654\ : std_logic;
signal \N__23647\ : std_logic;
signal \N__23646\ : std_logic;
signal \N__23645\ : std_logic;
signal \N__23642\ : std_logic;
signal \N__23639\ : std_logic;
signal \N__23638\ : std_logic;
signal \N__23637\ : std_logic;
signal \N__23634\ : std_logic;
signal \N__23631\ : std_logic;
signal \N__23628\ : std_logic;
signal \N__23623\ : std_logic;
signal \N__23614\ : std_logic;
signal \N__23611\ : std_logic;
signal \N__23608\ : std_logic;
signal \N__23605\ : std_logic;
signal \N__23602\ : std_logic;
signal \N__23599\ : std_logic;
signal \N__23596\ : std_logic;
signal \N__23595\ : std_logic;
signal \N__23592\ : std_logic;
signal \N__23589\ : std_logic;
signal \N__23586\ : std_logic;
signal \N__23581\ : std_logic;
signal \N__23578\ : std_logic;
signal \N__23575\ : std_logic;
signal \N__23572\ : std_logic;
signal \N__23571\ : std_logic;
signal \N__23566\ : std_logic;
signal \N__23563\ : std_logic;
signal \N__23560\ : std_logic;
signal \N__23557\ : std_logic;
signal \N__23554\ : std_logic;
signal \N__23551\ : std_logic;
signal \N__23550\ : std_logic;
signal \N__23549\ : std_logic;
signal \N__23542\ : std_logic;
signal \N__23539\ : std_logic;
signal \N__23536\ : std_logic;
signal \N__23533\ : std_logic;
signal \N__23530\ : std_logic;
signal \N__23527\ : std_logic;
signal \N__23524\ : std_logic;
signal \N__23521\ : std_logic;
signal \N__23518\ : std_logic;
signal \N__23515\ : std_logic;
signal \N__23512\ : std_logic;
signal \N__23509\ : std_logic;
signal \N__23506\ : std_logic;
signal \N__23503\ : std_logic;
signal \N__23500\ : std_logic;
signal \N__23497\ : std_logic;
signal \N__23494\ : std_logic;
signal \N__23491\ : std_logic;
signal \N__23488\ : std_logic;
signal \N__23485\ : std_logic;
signal \N__23482\ : std_logic;
signal \N__23479\ : std_logic;
signal \N__23478\ : std_logic;
signal \N__23477\ : std_logic;
signal \N__23476\ : std_logic;
signal \N__23473\ : std_logic;
signal \N__23470\ : std_logic;
signal \N__23465\ : std_logic;
signal \N__23458\ : std_logic;
signal \N__23457\ : std_logic;
signal \N__23456\ : std_logic;
signal \N__23455\ : std_logic;
signal \N__23454\ : std_logic;
signal \N__23453\ : std_logic;
signal \N__23452\ : std_logic;
signal \N__23449\ : std_logic;
signal \N__23448\ : std_logic;
signal \N__23447\ : std_logic;
signal \N__23446\ : std_logic;
signal \N__23445\ : std_logic;
signal \N__23444\ : std_logic;
signal \N__23441\ : std_logic;
signal \N__23440\ : std_logic;
signal \N__23439\ : std_logic;
signal \N__23438\ : std_logic;
signal \N__23437\ : std_logic;
signal \N__23436\ : std_logic;
signal \N__23435\ : std_logic;
signal \N__23432\ : std_logic;
signal \N__23431\ : std_logic;
signal \N__23430\ : std_logic;
signal \N__23423\ : std_logic;
signal \N__23422\ : std_logic;
signal \N__23415\ : std_logic;
signal \N__23412\ : std_logic;
signal \N__23405\ : std_logic;
signal \N__23402\ : std_logic;
signal \N__23397\ : std_logic;
signal \N__23390\ : std_logic;
signal \N__23389\ : std_logic;
signal \N__23388\ : std_logic;
signal \N__23385\ : std_logic;
signal \N__23382\ : std_logic;
signal \N__23381\ : std_logic;
signal \N__23378\ : std_logic;
signal \N__23377\ : std_logic;
signal \N__23376\ : std_logic;
signal \N__23375\ : std_logic;
signal \N__23372\ : std_logic;
signal \N__23369\ : std_logic;
signal \N__23366\ : std_logic;
signal \N__23363\ : std_logic;
signal \N__23358\ : std_logic;
signal \N__23351\ : std_logic;
signal \N__23346\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23344\ : std_logic;
signal \N__23343\ : std_logic;
signal \N__23342\ : std_logic;
signal \N__23341\ : std_logic;
signal \N__23340\ : std_logic;
signal \N__23337\ : std_logic;
signal \N__23334\ : std_logic;
signal \N__23331\ : std_logic;
signal \N__23328\ : std_logic;
signal \N__23327\ : std_logic;
signal \N__23326\ : std_logic;
signal \N__23321\ : std_logic;
signal \N__23318\ : std_logic;
signal \N__23315\ : std_logic;
signal \N__23308\ : std_logic;
signal \N__23301\ : std_logic;
signal \N__23298\ : std_logic;
signal \N__23295\ : std_logic;
signal \N__23286\ : std_logic;
signal \N__23277\ : std_logic;
signal \N__23272\ : std_logic;
signal \N__23261\ : std_logic;
signal \N__23248\ : std_logic;
signal \N__23247\ : std_logic;
signal \N__23246\ : std_logic;
signal \N__23241\ : std_logic;
signal \N__23240\ : std_logic;
signal \N__23239\ : std_logic;
signal \N__23236\ : std_logic;
signal \N__23235\ : std_logic;
signal \N__23234\ : std_logic;
signal \N__23233\ : std_logic;
signal \N__23232\ : std_logic;
signal \N__23229\ : std_logic;
signal \N__23224\ : std_logic;
signal \N__23223\ : std_logic;
signal \N__23222\ : std_logic;
signal \N__23221\ : std_logic;
signal \N__23220\ : std_logic;
signal \N__23217\ : std_logic;
signal \N__23214\ : std_logic;
signal \N__23207\ : std_logic;
signal \N__23202\ : std_logic;
signal \N__23199\ : std_logic;
signal \N__23192\ : std_logic;
signal \N__23187\ : std_logic;
signal \N__23176\ : std_logic;
signal \N__23175\ : std_logic;
signal \N__23174\ : std_logic;
signal \N__23171\ : std_logic;
signal \N__23170\ : std_logic;
signal \N__23163\ : std_logic;
signal \N__23162\ : std_logic;
signal \N__23161\ : std_logic;
signal \N__23158\ : std_logic;
signal \N__23157\ : std_logic;
signal \N__23154\ : std_logic;
signal \N__23147\ : std_logic;
signal \N__23144\ : std_logic;
signal \N__23141\ : std_logic;
signal \N__23138\ : std_logic;
signal \N__23131\ : std_logic;
signal \N__23130\ : std_logic;
signal \N__23127\ : std_logic;
signal \N__23124\ : std_logic;
signal \N__23121\ : std_logic;
signal \N__23118\ : std_logic;
signal \N__23113\ : std_logic;
signal \N__23112\ : std_logic;
signal \N__23109\ : std_logic;
signal \N__23106\ : std_logic;
signal \N__23105\ : std_logic;
signal \N__23102\ : std_logic;
signal \N__23097\ : std_logic;
signal \N__23092\ : std_logic;
signal \N__23091\ : std_logic;
signal \N__23090\ : std_logic;
signal \N__23087\ : std_logic;
signal \N__23082\ : std_logic;
signal \N__23077\ : std_logic;
signal \N__23076\ : std_logic;
signal \N__23075\ : std_logic;
signal \N__23072\ : std_logic;
signal \N__23069\ : std_logic;
signal \N__23066\ : std_logic;
signal \N__23059\ : std_logic;
signal \N__23058\ : std_logic;
signal \N__23057\ : std_logic;
signal \N__23054\ : std_logic;
signal \N__23051\ : std_logic;
signal \N__23048\ : std_logic;
signal \N__23045\ : std_logic;
signal \N__23038\ : std_logic;
signal \N__23037\ : std_logic;
signal \N__23036\ : std_logic;
signal \N__23033\ : std_logic;
signal \N__23030\ : std_logic;
signal \N__23027\ : std_logic;
signal \N__23020\ : std_logic;
signal \N__23019\ : std_logic;
signal \N__23018\ : std_logic;
signal \N__23015\ : std_logic;
signal \N__23014\ : std_logic;
signal \N__23011\ : std_logic;
signal \N__23008\ : std_logic;
signal \N__23003\ : std_logic;
signal \N__22998\ : std_logic;
signal \N__22995\ : std_logic;
signal \N__22992\ : std_logic;
signal \N__22989\ : std_logic;
signal \N__22984\ : std_logic;
signal \N__22983\ : std_logic;
signal \N__22980\ : std_logic;
signal \N__22979\ : std_logic;
signal \N__22976\ : std_logic;
signal \N__22973\ : std_logic;
signal \N__22970\ : std_logic;
signal \N__22963\ : std_logic;
signal \N__22962\ : std_logic;
signal \N__22961\ : std_logic;
signal \N__22954\ : std_logic;
signal \N__22953\ : std_logic;
signal \N__22950\ : std_logic;
signal \N__22947\ : std_logic;
signal \N__22944\ : std_logic;
signal \N__22941\ : std_logic;
signal \N__22938\ : std_logic;
signal \N__22935\ : std_logic;
signal \N__22930\ : std_logic;
signal \N__22929\ : std_logic;
signal \N__22926\ : std_logic;
signal \N__22925\ : std_logic;
signal \N__22922\ : std_logic;
signal \N__22919\ : std_logic;
signal \N__22916\ : std_logic;
signal \N__22909\ : std_logic;
signal \N__22908\ : std_logic;
signal \N__22907\ : std_logic;
signal \N__22906\ : std_logic;
signal \N__22897\ : std_logic;
signal \N__22894\ : std_logic;
signal \N__22891\ : std_logic;
signal \N__22888\ : std_logic;
signal \N__22885\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22881\ : std_logic;
signal \N__22878\ : std_logic;
signal \N__22875\ : std_logic;
signal \N__22874\ : std_logic;
signal \N__22873\ : std_logic;
signal \N__22864\ : std_logic;
signal \N__22861\ : std_logic;
signal \N__22858\ : std_logic;
signal \N__22855\ : std_logic;
signal \N__22854\ : std_logic;
signal \N__22851\ : std_logic;
signal \N__22848\ : std_logic;
signal \N__22843\ : std_logic;
signal \N__22840\ : std_logic;
signal \N__22837\ : std_logic;
signal \N__22834\ : std_logic;
signal \N__22831\ : std_logic;
signal \N__22828\ : std_logic;
signal \N__22827\ : std_logic;
signal \N__22824\ : std_logic;
signal \N__22821\ : std_logic;
signal \N__22820\ : std_logic;
signal \N__22815\ : std_logic;
signal \N__22812\ : std_logic;
signal \N__22807\ : std_logic;
signal \N__22806\ : std_logic;
signal \N__22803\ : std_logic;
signal \N__22800\ : std_logic;
signal \N__22797\ : std_logic;
signal \N__22794\ : std_logic;
signal \N__22793\ : std_logic;
signal \N__22792\ : std_logic;
signal \N__22787\ : std_logic;
signal \N__22784\ : std_logic;
signal \N__22781\ : std_logic;
signal \N__22776\ : std_logic;
signal \N__22773\ : std_logic;
signal \N__22770\ : std_logic;
signal \N__22765\ : std_logic;
signal \N__22764\ : std_logic;
signal \N__22761\ : std_logic;
signal \N__22760\ : std_logic;
signal \N__22757\ : std_logic;
signal \N__22754\ : std_logic;
signal \N__22751\ : std_logic;
signal \N__22748\ : std_logic;
signal \N__22745\ : std_logic;
signal \N__22738\ : std_logic;
signal \N__22735\ : std_logic;
signal \N__22734\ : std_logic;
signal \N__22733\ : std_logic;
signal \N__22730\ : std_logic;
signal \N__22727\ : std_logic;
signal \N__22724\ : std_logic;
signal \N__22721\ : std_logic;
signal \N__22714\ : std_logic;
signal \N__22713\ : std_logic;
signal \N__22712\ : std_logic;
signal \N__22711\ : std_logic;
signal \N__22702\ : std_logic;
signal \N__22699\ : std_logic;
signal \N__22696\ : std_logic;
signal \N__22693\ : std_logic;
signal \N__22690\ : std_logic;
signal \N__22689\ : std_logic;
signal \N__22688\ : std_logic;
signal \N__22685\ : std_logic;
signal \N__22682\ : std_logic;
signal \N__22679\ : std_logic;
signal \N__22676\ : std_logic;
signal \N__22669\ : std_logic;
signal \N__22666\ : std_logic;
signal \N__22665\ : std_logic;
signal \N__22662\ : std_logic;
signal \N__22661\ : std_logic;
signal \N__22658\ : std_logic;
signal \N__22655\ : std_logic;
signal \N__22652\ : std_logic;
signal \N__22649\ : std_logic;
signal \N__22642\ : std_logic;
signal \N__22639\ : std_logic;
signal \N__22636\ : std_logic;
signal \N__22633\ : std_logic;
signal \N__22632\ : std_logic;
signal \N__22631\ : std_logic;
signal \N__22628\ : std_logic;
signal \N__22623\ : std_logic;
signal \N__22618\ : std_logic;
signal \N__22615\ : std_logic;
signal \N__22614\ : std_logic;
signal \N__22613\ : std_logic;
signal \N__22610\ : std_logic;
signal \N__22605\ : std_logic;
signal \N__22600\ : std_logic;
signal \N__22597\ : std_logic;
signal \N__22596\ : std_logic;
signal \N__22595\ : std_logic;
signal \N__22594\ : std_logic;
signal \N__22593\ : std_logic;
signal \N__22582\ : std_logic;
signal \N__22579\ : std_logic;
signal \N__22578\ : std_logic;
signal \N__22577\ : std_logic;
signal \N__22576\ : std_logic;
signal \N__22569\ : std_logic;
signal \N__22566\ : std_logic;
signal \N__22561\ : std_logic;
signal \N__22560\ : std_logic;
signal \N__22557\ : std_logic;
signal \N__22556\ : std_logic;
signal \N__22551\ : std_logic;
signal \N__22548\ : std_logic;
signal \N__22543\ : std_logic;
signal \N__22540\ : std_logic;
signal \N__22539\ : std_logic;
signal \N__22538\ : std_logic;
signal \N__22537\ : std_logic;
signal \N__22534\ : std_logic;
signal \N__22525\ : std_logic;
signal \N__22522\ : std_logic;
signal \N__22521\ : std_logic;
signal \N__22520\ : std_logic;
signal \N__22519\ : std_logic;
signal \N__22516\ : std_logic;
signal \N__22515\ : std_logic;
signal \N__22506\ : std_logic;
signal \N__22503\ : std_logic;
signal \N__22498\ : std_logic;
signal \N__22495\ : std_logic;
signal \N__22492\ : std_logic;
signal \N__22489\ : std_logic;
signal \N__22488\ : std_logic;
signal \N__22487\ : std_logic;
signal \N__22486\ : std_logic;
signal \N__22481\ : std_logic;
signal \N__22478\ : std_logic;
signal \N__22475\ : std_logic;
signal \N__22472\ : std_logic;
signal \N__22469\ : std_logic;
signal \N__22462\ : std_logic;
signal \N__22461\ : std_logic;
signal \N__22460\ : std_logic;
signal \N__22459\ : std_logic;
signal \N__22456\ : std_logic;
signal \N__22455\ : std_logic;
signal \N__22450\ : std_logic;
signal \N__22447\ : std_logic;
signal \N__22442\ : std_logic;
signal \N__22439\ : std_logic;
signal \N__22436\ : std_logic;
signal \N__22429\ : std_logic;
signal \N__22428\ : std_logic;
signal \N__22427\ : std_logic;
signal \N__22426\ : std_logic;
signal \N__22425\ : std_logic;
signal \N__22424\ : std_logic;
signal \N__22423\ : std_logic;
signal \N__22416\ : std_logic;
signal \N__22409\ : std_logic;
signal \N__22406\ : std_logic;
signal \N__22399\ : std_logic;
signal \N__22398\ : std_logic;
signal \N__22397\ : std_logic;
signal \N__22396\ : std_logic;
signal \N__22395\ : std_logic;
signal \N__22390\ : std_logic;
signal \N__22383\ : std_logic;
signal \N__22378\ : std_logic;
signal \N__22375\ : std_logic;
signal \N__22374\ : std_logic;
signal \N__22371\ : std_logic;
signal \N__22370\ : std_logic;
signal \N__22367\ : std_logic;
signal \N__22364\ : std_logic;
signal \N__22359\ : std_logic;
signal \N__22354\ : std_logic;
signal \N__22353\ : std_logic;
signal \N__22352\ : std_logic;
signal \N__22351\ : std_logic;
signal \N__22350\ : std_logic;
signal \N__22343\ : std_logic;
signal \N__22340\ : std_logic;
signal \N__22337\ : std_logic;
signal \N__22332\ : std_logic;
signal \N__22327\ : std_logic;
signal \N__22326\ : std_logic;
signal \N__22323\ : std_logic;
signal \N__22322\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22313\ : std_logic;
signal \N__22312\ : std_logic;
signal \N__22307\ : std_logic;
signal \N__22304\ : std_logic;
signal \N__22301\ : std_logic;
signal \N__22294\ : std_logic;
signal \N__22293\ : std_logic;
signal \N__22292\ : std_logic;
signal \N__22285\ : std_logic;
signal \N__22282\ : std_logic;
signal \N__22281\ : std_logic;
signal \N__22280\ : std_logic;
signal \N__22277\ : std_logic;
signal \N__22272\ : std_logic;
signal \N__22269\ : std_logic;
signal \N__22264\ : std_logic;
signal \N__22261\ : std_logic;
signal \N__22260\ : std_logic;
signal \N__22259\ : std_logic;
signal \N__22256\ : std_logic;
signal \N__22251\ : std_logic;
signal \N__22248\ : std_logic;
signal \N__22243\ : std_logic;
signal \N__22242\ : std_logic;
signal \N__22241\ : std_logic;
signal \N__22236\ : std_logic;
signal \N__22235\ : std_logic;
signal \N__22232\ : std_logic;
signal \N__22229\ : std_logic;
signal \N__22226\ : std_logic;
signal \N__22219\ : std_logic;
signal \N__22216\ : std_logic;
signal \N__22215\ : std_logic;
signal \N__22214\ : std_logic;
signal \N__22213\ : std_logic;
signal \N__22208\ : std_logic;
signal \N__22205\ : std_logic;
signal \N__22202\ : std_logic;
signal \N__22195\ : std_logic;
signal \N__22194\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22192\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22184\ : std_logic;
signal \N__22181\ : std_logic;
signal \N__22174\ : std_logic;
signal \N__22173\ : std_logic;
signal \N__22172\ : std_logic;
signal \N__22171\ : std_logic;
signal \N__22170\ : std_logic;
signal \N__22159\ : std_logic;
signal \N__22156\ : std_logic;
signal \N__22153\ : std_logic;
signal \N__22150\ : std_logic;
signal \N__22147\ : std_logic;
signal \N__22146\ : std_logic;
signal \N__22143\ : std_logic;
signal \N__22140\ : std_logic;
signal \N__22135\ : std_logic;
signal \N__22132\ : std_logic;
signal \N__22129\ : std_logic;
signal \N__22128\ : std_logic;
signal \N__22127\ : std_logic;
signal \N__22124\ : std_logic;
signal \N__22121\ : std_logic;
signal \N__22118\ : std_logic;
signal \N__22111\ : std_logic;
signal \N__22110\ : std_logic;
signal \N__22109\ : std_logic;
signal \N__22106\ : std_logic;
signal \N__22103\ : std_logic;
signal \N__22096\ : std_logic;
signal \N__22093\ : std_logic;
signal \N__22092\ : std_logic;
signal \N__22091\ : std_logic;
signal \N__22090\ : std_logic;
signal \N__22083\ : std_logic;
signal \N__22080\ : std_logic;
signal \N__22075\ : std_logic;
signal \N__22072\ : std_logic;
signal \N__22071\ : std_logic;
signal \N__22068\ : std_logic;
signal \N__22065\ : std_logic;
signal \N__22062\ : std_logic;
signal \N__22057\ : std_logic;
signal \N__22056\ : std_logic;
signal \N__22055\ : std_logic;
signal \N__22052\ : std_logic;
signal \N__22049\ : std_logic;
signal \N__22046\ : std_logic;
signal \N__22039\ : std_logic;
signal \N__22036\ : std_logic;
signal \N__22035\ : std_logic;
signal \N__22034\ : std_logic;
signal \N__22033\ : std_logic;
signal \N__22026\ : std_logic;
signal \N__22023\ : std_logic;
signal \N__22018\ : std_logic;
signal \N__22015\ : std_logic;
signal \N__22012\ : std_logic;
signal \N__22009\ : std_logic;
signal \N__22006\ : std_logic;
signal \N__22003\ : std_logic;
signal \N__22000\ : std_logic;
signal \N__21999\ : std_logic;
signal \N__21996\ : std_logic;
signal \N__21995\ : std_logic;
signal \N__21992\ : std_logic;
signal \N__21991\ : std_logic;
signal \N__21988\ : std_logic;
signal \N__21987\ : std_logic;
signal \N__21986\ : std_logic;
signal \N__21983\ : std_logic;
signal \N__21980\ : std_logic;
signal \N__21977\ : std_logic;
signal \N__21974\ : std_logic;
signal \N__21971\ : std_logic;
signal \N__21966\ : std_logic;
signal \N__21963\ : std_logic;
signal \N__21960\ : std_logic;
signal \N__21957\ : std_logic;
signal \N__21954\ : std_logic;
signal \N__21949\ : std_logic;
signal \N__21946\ : std_logic;
signal \N__21937\ : std_logic;
signal \N__21936\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21932\ : std_logic;
signal \N__21929\ : std_logic;
signal \N__21926\ : std_logic;
signal \N__21925\ : std_logic;
signal \N__21924\ : std_logic;
signal \N__21919\ : std_logic;
signal \N__21918\ : std_logic;
signal \N__21915\ : std_logic;
signal \N__21910\ : std_logic;
signal \N__21907\ : std_logic;
signal \N__21904\ : std_logic;
signal \N__21895\ : std_logic;
signal \N__21892\ : std_logic;
signal \N__21891\ : std_logic;
signal \N__21888\ : std_logic;
signal \N__21885\ : std_logic;
signal \N__21882\ : std_logic;
signal \N__21877\ : std_logic;
signal \N__21876\ : std_logic;
signal \N__21873\ : std_logic;
signal \N__21872\ : std_logic;
signal \N__21871\ : std_logic;
signal \N__21868\ : std_logic;
signal \N__21865\ : std_logic;
signal \N__21862\ : std_logic;
signal \N__21859\ : std_logic;
signal \N__21852\ : std_logic;
signal \N__21849\ : std_logic;
signal \N__21846\ : std_logic;
signal \N__21841\ : std_logic;
signal \N__21838\ : std_logic;
signal \N__21837\ : std_logic;
signal \N__21834\ : std_logic;
signal \N__21833\ : std_logic;
signal \N__21832\ : std_logic;
signal \N__21831\ : std_logic;
signal \N__21828\ : std_logic;
signal \N__21825\ : std_logic;
signal \N__21820\ : std_logic;
signal \N__21819\ : std_logic;
signal \N__21816\ : std_logic;
signal \N__21813\ : std_logic;
signal \N__21810\ : std_logic;
signal \N__21807\ : std_logic;
signal \N__21802\ : std_logic;
signal \N__21793\ : std_logic;
signal \N__21790\ : std_logic;
signal \N__21787\ : std_logic;
signal \N__21784\ : std_logic;
signal \N__21781\ : std_logic;
signal \N__21780\ : std_logic;
signal \N__21777\ : std_logic;
signal \N__21774\ : std_logic;
signal \N__21771\ : std_logic;
signal \N__21768\ : std_logic;
signal \N__21767\ : std_logic;
signal \N__21766\ : std_logic;
signal \N__21765\ : std_logic;
signal \N__21764\ : std_logic;
signal \N__21763\ : std_logic;
signal \N__21760\ : std_logic;
signal \N__21757\ : std_logic;
signal \N__21756\ : std_logic;
signal \N__21753\ : std_logic;
signal \N__21750\ : std_logic;
signal \N__21749\ : std_logic;
signal \N__21742\ : std_logic;
signal \N__21739\ : std_logic;
signal \N__21736\ : std_logic;
signal \N__21727\ : std_logic;
signal \N__21718\ : std_logic;
signal \N__21715\ : std_logic;
signal \N__21712\ : std_logic;
signal \N__21709\ : std_logic;
signal \N__21706\ : std_logic;
signal \N__21703\ : std_logic;
signal \N__21700\ : std_logic;
signal \N__21699\ : std_logic;
signal \N__21698\ : std_logic;
signal \N__21697\ : std_logic;
signal \N__21696\ : std_logic;
signal \N__21695\ : std_logic;
signal \N__21692\ : std_logic;
signal \N__21689\ : std_logic;
signal \N__21686\ : std_logic;
signal \N__21685\ : std_logic;
signal \N__21684\ : std_logic;
signal \N__21683\ : std_logic;
signal \N__21680\ : std_logic;
signal \N__21675\ : std_logic;
signal \N__21672\ : std_logic;
signal \N__21669\ : std_logic;
signal \N__21660\ : std_logic;
signal \N__21649\ : std_logic;
signal \N__21646\ : std_logic;
signal \N__21643\ : std_logic;
signal \N__21640\ : std_logic;
signal \N__21637\ : std_logic;
signal \N__21634\ : std_logic;
signal \N__21631\ : std_logic;
signal \N__21628\ : std_logic;
signal \N__21625\ : std_logic;
signal \N__21624\ : std_logic;
signal \N__21623\ : std_logic;
signal \N__21622\ : std_logic;
signal \N__21621\ : std_logic;
signal \N__21620\ : std_logic;
signal \N__21619\ : std_logic;
signal \N__21618\ : std_logic;
signal \N__21617\ : std_logic;
signal \N__21616\ : std_logic;
signal \N__21615\ : std_logic;
signal \N__21614\ : std_logic;
signal \N__21611\ : std_logic;
signal \N__21610\ : std_logic;
signal \N__21609\ : std_logic;
signal \N__21608\ : std_logic;
signal \N__21607\ : std_logic;
signal \N__21606\ : std_logic;
signal \N__21603\ : std_logic;
signal \N__21598\ : std_logic;
signal \N__21581\ : std_logic;
signal \N__21578\ : std_logic;
signal \N__21577\ : std_logic;
signal \N__21576\ : std_logic;
signal \N__21575\ : std_logic;
signal \N__21574\ : std_logic;
signal \N__21573\ : std_logic;
signal \N__21572\ : std_logic;
signal \N__21569\ : std_logic;
signal \N__21568\ : std_logic;
signal \N__21565\ : std_logic;
signal \N__21562\ : std_logic;
signal \N__21559\ : std_logic;
signal \N__21556\ : std_logic;
signal \N__21553\ : std_logic;
signal \N__21550\ : std_logic;
signal \N__21547\ : std_logic;
signal \N__21544\ : std_logic;
signal \N__21537\ : std_logic;
signal \N__21536\ : std_logic;
signal \N__21529\ : std_logic;
signal \N__21522\ : std_logic;
signal \N__21521\ : std_logic;
signal \N__21520\ : std_logic;
signal \N__21519\ : std_logic;
signal \N__21518\ : std_logic;
signal \N__21517\ : std_logic;
signal \N__21516\ : std_logic;
signal \N__21515\ : std_logic;
signal \N__21514\ : std_logic;
signal \N__21513\ : std_logic;
signal \N__21508\ : std_logic;
signal \N__21501\ : std_logic;
signal \N__21496\ : std_logic;
signal \N__21493\ : std_logic;
signal \N__21490\ : std_logic;
signal \N__21485\ : std_logic;
signal \N__21470\ : std_logic;
signal \N__21465\ : std_logic;
signal \N__21462\ : std_logic;
signal \N__21445\ : std_logic;
signal \N__21444\ : std_logic;
signal \N__21443\ : std_logic;
signal \N__21442\ : std_logic;
signal \N__21441\ : std_logic;
signal \N__21438\ : std_logic;
signal \N__21435\ : std_logic;
signal \N__21430\ : std_logic;
signal \N__21427\ : std_logic;
signal \N__21420\ : std_logic;
signal \N__21415\ : std_logic;
signal \N__21414\ : std_logic;
signal \N__21411\ : std_logic;
signal \N__21408\ : std_logic;
signal \N__21407\ : std_logic;
signal \N__21406\ : std_logic;
signal \N__21403\ : std_logic;
signal \N__21400\ : std_logic;
signal \N__21395\ : std_logic;
signal \N__21394\ : std_logic;
signal \N__21393\ : std_logic;
signal \N__21392\ : std_logic;
signal \N__21391\ : std_logic;
signal \N__21390\ : std_logic;
signal \N__21389\ : std_logic;
signal \N__21384\ : std_logic;
signal \N__21381\ : std_logic;
signal \N__21376\ : std_logic;
signal \N__21367\ : std_logic;
signal \N__21358\ : std_logic;
signal \N__21355\ : std_logic;
signal \N__21352\ : std_logic;
signal \N__21351\ : std_logic;
signal \N__21348\ : std_logic;
signal \N__21347\ : std_logic;
signal \N__21346\ : std_logic;
signal \N__21343\ : std_logic;
signal \N__21340\ : std_logic;
signal \N__21335\ : std_logic;
signal \N__21330\ : std_logic;
signal \N__21325\ : std_logic;
signal \N__21322\ : std_logic;
signal \N__21319\ : std_logic;
signal \N__21316\ : std_logic;
signal \N__21313\ : std_logic;
signal \N__21310\ : std_logic;
signal \N__21307\ : std_logic;
signal \N__21304\ : std_logic;
signal \N__21301\ : std_logic;
signal \N__21298\ : std_logic;
signal \N__21295\ : std_logic;
signal \N__21292\ : std_logic;
signal \N__21291\ : std_logic;
signal \N__21290\ : std_logic;
signal \N__21287\ : std_logic;
signal \N__21286\ : std_logic;
signal \N__21281\ : std_logic;
signal \N__21278\ : std_logic;
signal \N__21275\ : std_logic;
signal \N__21268\ : std_logic;
signal \N__21267\ : std_logic;
signal \N__21266\ : std_logic;
signal \N__21265\ : std_logic;
signal \N__21264\ : std_logic;
signal \N__21261\ : std_logic;
signal \N__21260\ : std_logic;
signal \N__21259\ : std_logic;
signal \N__21254\ : std_logic;
signal \N__21251\ : std_logic;
signal \N__21250\ : std_logic;
signal \N__21247\ : std_logic;
signal \N__21246\ : std_logic;
signal \N__21245\ : std_logic;
signal \N__21244\ : std_logic;
signal \N__21241\ : std_logic;
signal \N__21238\ : std_logic;
signal \N__21235\ : std_logic;
signal \N__21234\ : std_logic;
signal \N__21231\ : std_logic;
signal \N__21228\ : std_logic;
signal \N__21223\ : std_logic;
signal \N__21222\ : std_logic;
signal \N__21219\ : std_logic;
signal \N__21218\ : std_logic;
signal \N__21215\ : std_logic;
signal \N__21212\ : std_logic;
signal \N__21207\ : std_logic;
signal \N__21204\ : std_logic;
signal \N__21201\ : std_logic;
signal \N__21194\ : std_logic;
signal \N__21191\ : std_logic;
signal \N__21188\ : std_logic;
signal \N__21185\ : std_logic;
signal \N__21182\ : std_logic;
signal \N__21179\ : std_logic;
signal \N__21176\ : std_logic;
signal \N__21171\ : std_logic;
signal \N__21168\ : std_logic;
signal \N__21165\ : std_logic;
signal \N__21160\ : std_logic;
signal \N__21157\ : std_logic;
signal \N__21152\ : std_logic;
signal \N__21147\ : std_logic;
signal \N__21136\ : std_logic;
signal \N__21133\ : std_logic;
signal \N__21130\ : std_logic;
signal \N__21127\ : std_logic;
signal \N__21124\ : std_logic;
signal \N__21121\ : std_logic;
signal \N__21118\ : std_logic;
signal \N__21115\ : std_logic;
signal \N__21112\ : std_logic;
signal \N__21111\ : std_logic;
signal \N__21110\ : std_logic;
signal \N__21109\ : std_logic;
signal \N__21108\ : std_logic;
signal \N__21107\ : std_logic;
signal \N__21104\ : std_logic;
signal \N__21099\ : std_logic;
signal \N__21098\ : std_logic;
signal \N__21097\ : std_logic;
signal \N__21096\ : std_logic;
signal \N__21095\ : std_logic;
signal \N__21094\ : std_logic;
signal \N__21093\ : std_logic;
signal \N__21092\ : std_logic;
signal \N__21091\ : std_logic;
signal \N__21090\ : std_logic;
signal \N__21087\ : std_logic;
signal \N__21084\ : std_logic;
signal \N__21081\ : std_logic;
signal \N__21076\ : std_logic;
signal \N__21073\ : std_logic;
signal \N__21072\ : std_logic;
signal \N__21071\ : std_logic;
signal \N__21054\ : std_logic;
signal \N__21051\ : std_logic;
signal \N__21048\ : std_logic;
signal \N__21045\ : std_logic;
signal \N__21044\ : std_logic;
signal \N__21043\ : std_logic;
signal \N__21042\ : std_logic;
signal \N__21041\ : std_logic;
signal \N__21040\ : std_logic;
signal \N__21039\ : std_logic;
signal \N__21038\ : std_logic;
signal \N__21037\ : std_logic;
signal \N__21036\ : std_logic;
signal \N__21035\ : std_logic;
signal \N__21034\ : std_logic;
signal \N__21033\ : std_logic;
signal \N__21032\ : std_logic;
signal \N__21031\ : std_logic;
signal \N__21030\ : std_logic;
signal \N__21029\ : std_logic;
signal \N__21028\ : std_logic;
signal \N__21023\ : std_logic;
signal \N__21020\ : std_logic;
signal \N__21017\ : std_logic;
signal \N__21008\ : std_logic;
signal \N__21001\ : std_logic;
signal \N__20990\ : std_logic;
signal \N__20985\ : std_logic;
signal \N__20970\ : std_logic;
signal \N__20967\ : std_logic;
signal \N__20950\ : std_logic;
signal \N__20949\ : std_logic;
signal \N__20946\ : std_logic;
signal \N__20941\ : std_logic;
signal \N__20940\ : std_logic;
signal \N__20939\ : std_logic;
signal \N__20938\ : std_logic;
signal \N__20937\ : std_logic;
signal \N__20936\ : std_logic;
signal \N__20935\ : std_logic;
signal \N__20932\ : std_logic;
signal \N__20929\ : std_logic;
signal \N__20926\ : std_logic;
signal \N__20923\ : std_logic;
signal \N__20916\ : std_logic;
signal \N__20913\ : std_logic;
signal \N__20910\ : std_logic;
signal \N__20907\ : std_logic;
signal \N__20904\ : std_logic;
signal \N__20901\ : std_logic;
signal \N__20900\ : std_logic;
signal \N__20895\ : std_logic;
signal \N__20892\ : std_logic;
signal \N__20891\ : std_logic;
signal \N__20886\ : std_logic;
signal \N__20883\ : std_logic;
signal \N__20880\ : std_logic;
signal \N__20877\ : std_logic;
signal \N__20874\ : std_logic;
signal \N__20871\ : std_logic;
signal \N__20860\ : std_logic;
signal \N__20857\ : std_logic;
signal \N__20854\ : std_logic;
signal \N__20851\ : std_logic;
signal \N__20848\ : std_logic;
signal \N__20845\ : std_logic;
signal \N__20842\ : std_logic;
signal \N__20839\ : std_logic;
signal \N__20838\ : std_logic;
signal \N__20835\ : std_logic;
signal \N__20832\ : std_logic;
signal \N__20829\ : std_logic;
signal \N__20824\ : std_logic;
signal \N__20821\ : std_logic;
signal \N__20818\ : std_logic;
signal \N__20815\ : std_logic;
signal \N__20814\ : std_logic;
signal \N__20813\ : std_logic;
signal \N__20812\ : std_logic;
signal \N__20811\ : std_logic;
signal \N__20810\ : std_logic;
signal \N__20809\ : std_logic;
signal \N__20808\ : std_logic;
signal \N__20807\ : std_logic;
signal \N__20806\ : std_logic;
signal \N__20805\ : std_logic;
signal \N__20802\ : std_logic;
signal \N__20799\ : std_logic;
signal \N__20796\ : std_logic;
signal \N__20795\ : std_logic;
signal \N__20794\ : std_logic;
signal \N__20793\ : std_logic;
signal \N__20792\ : std_logic;
signal \N__20789\ : std_logic;
signal \N__20786\ : std_logic;
signal \N__20783\ : std_logic;
signal \N__20780\ : std_logic;
signal \N__20777\ : std_logic;
signal \N__20774\ : std_logic;
signal \N__20771\ : std_logic;
signal \N__20768\ : std_logic;
signal \N__20767\ : std_logic;
signal \N__20764\ : std_logic;
signal \N__20761\ : std_logic;
signal \N__20758\ : std_logic;
signal \N__20757\ : std_logic;
signal \N__20756\ : std_logic;
signal \N__20755\ : std_logic;
signal \N__20752\ : std_logic;
signal \N__20751\ : std_logic;
signal \N__20748\ : std_logic;
signal \N__20747\ : std_logic;
signal \N__20746\ : std_logic;
signal \N__20743\ : std_logic;
signal \N__20742\ : std_logic;
signal \N__20739\ : std_logic;
signal \N__20730\ : std_logic;
signal \N__20721\ : std_logic;
signal \N__20718\ : std_logic;
signal \N__20713\ : std_logic;
signal \N__20710\ : std_logic;
signal \N__20705\ : std_logic;
signal \N__20698\ : std_logic;
signal \N__20685\ : std_logic;
signal \N__20668\ : std_logic;
signal \N__20667\ : std_logic;
signal \N__20666\ : std_logic;
signal \N__20665\ : std_logic;
signal \N__20664\ : std_logic;
signal \N__20663\ : std_logic;
signal \N__20662\ : std_logic;
signal \N__20661\ : std_logic;
signal \N__20660\ : std_logic;
signal \N__20659\ : std_logic;
signal \N__20658\ : std_logic;
signal \N__20657\ : std_logic;
signal \N__20654\ : std_logic;
signal \N__20653\ : std_logic;
signal \N__20644\ : std_logic;
signal \N__20635\ : std_logic;
signal \N__20634\ : std_logic;
signal \N__20631\ : std_logic;
signal \N__20628\ : std_logic;
signal \N__20627\ : std_logic;
signal \N__20624\ : std_logic;
signal \N__20623\ : std_logic;
signal \N__20622\ : std_logic;
signal \N__20619\ : std_logic;
signal \N__20616\ : std_logic;
signal \N__20611\ : std_logic;
signal \N__20598\ : std_logic;
signal \N__20595\ : std_logic;
signal \N__20592\ : std_logic;
signal \N__20585\ : std_logic;
signal \N__20578\ : std_logic;
signal \N__20575\ : std_logic;
signal \N__20572\ : std_logic;
signal \N__20569\ : std_logic;
signal \N__20566\ : std_logic;
signal \N__20563\ : std_logic;
signal \N__20562\ : std_logic;
signal \N__20561\ : std_logic;
signal \N__20560\ : std_logic;
signal \N__20557\ : std_logic;
signal \N__20554\ : std_logic;
signal \N__20551\ : std_logic;
signal \N__20548\ : std_logic;
signal \N__20539\ : std_logic;
signal \N__20536\ : std_logic;
signal \N__20533\ : std_logic;
signal \N__20530\ : std_logic;
signal \N__20529\ : std_logic;
signal \N__20524\ : std_logic;
signal \N__20521\ : std_logic;
signal \N__20518\ : std_logic;
signal \N__20517\ : std_logic;
signal \N__20516\ : std_logic;
signal \N__20515\ : std_logic;
signal \N__20508\ : std_logic;
signal \N__20507\ : std_logic;
signal \N__20506\ : std_logic;
signal \N__20503\ : std_logic;
signal \N__20500\ : std_logic;
signal \N__20495\ : std_logic;
signal \N__20492\ : std_logic;
signal \N__20487\ : std_logic;
signal \N__20484\ : std_logic;
signal \N__20481\ : std_logic;
signal \N__20476\ : std_logic;
signal \N__20475\ : std_logic;
signal \N__20472\ : std_logic;
signal \N__20469\ : std_logic;
signal \N__20466\ : std_logic;
signal \N__20463\ : std_logic;
signal \N__20458\ : std_logic;
signal \N__20457\ : std_logic;
signal \N__20454\ : std_logic;
signal \N__20451\ : std_logic;
signal \N__20448\ : std_logic;
signal \N__20445\ : std_logic;
signal \N__20442\ : std_logic;
signal \N__20437\ : std_logic;
signal \N__20434\ : std_logic;
signal \N__20433\ : std_logic;
signal \N__20428\ : std_logic;
signal \N__20425\ : std_logic;
signal \N__20424\ : std_logic;
signal \N__20423\ : std_logic;
signal \N__20422\ : std_logic;
signal \N__20419\ : std_logic;
signal \N__20412\ : std_logic;
signal \N__20409\ : std_logic;
signal \N__20406\ : std_logic;
signal \N__20401\ : std_logic;
signal \N__20398\ : std_logic;
signal \N__20397\ : std_logic;
signal \N__20396\ : std_logic;
signal \N__20395\ : std_logic;
signal \N__20394\ : std_logic;
signal \N__20393\ : std_logic;
signal \N__20392\ : std_logic;
signal \N__20389\ : std_logic;
signal \N__20388\ : std_logic;
signal \N__20385\ : std_logic;
signal \N__20382\ : std_logic;
signal \N__20379\ : std_logic;
signal \N__20374\ : std_logic;
signal \N__20371\ : std_logic;
signal \N__20370\ : std_logic;
signal \N__20369\ : std_logic;
signal \N__20362\ : std_logic;
signal \N__20361\ : std_logic;
signal \N__20360\ : std_logic;
signal \N__20357\ : std_logic;
signal \N__20352\ : std_logic;
signal \N__20349\ : std_logic;
signal \N__20346\ : std_logic;
signal \N__20343\ : std_logic;
signal \N__20340\ : std_logic;
signal \N__20335\ : std_logic;
signal \N__20334\ : std_logic;
signal \N__20329\ : std_logic;
signal \N__20324\ : std_logic;
signal \N__20321\ : std_logic;
signal \N__20316\ : std_logic;
signal \N__20313\ : std_logic;
signal \N__20308\ : std_logic;
signal \N__20299\ : std_logic;
signal \N__20296\ : std_logic;
signal \N__20295\ : std_logic;
signal \N__20292\ : std_logic;
signal \N__20289\ : std_logic;
signal \N__20284\ : std_logic;
signal \N__20283\ : std_logic;
signal \N__20280\ : std_logic;
signal \N__20277\ : std_logic;
signal \N__20274\ : std_logic;
signal \N__20271\ : std_logic;
signal \N__20268\ : std_logic;
signal \N__20263\ : std_logic;
signal \N__20260\ : std_logic;
signal \N__20257\ : std_logic;
signal \N__20254\ : std_logic;
signal \N__20251\ : std_logic;
signal \N__20248\ : std_logic;
signal \N__20245\ : std_logic;
signal \N__20242\ : std_logic;
signal \N__20239\ : std_logic;
signal \N__20236\ : std_logic;
signal \N__20235\ : std_logic;
signal \N__20230\ : std_logic;
signal \N__20227\ : std_logic;
signal \N__20224\ : std_logic;
signal \N__20223\ : std_logic;
signal \N__20220\ : std_logic;
signal \N__20217\ : std_logic;
signal \N__20212\ : std_logic;
signal \N__20209\ : std_logic;
signal \N__20206\ : std_logic;
signal \N__20203\ : std_logic;
signal \N__20200\ : std_logic;
signal \N__20197\ : std_logic;
signal \N__20194\ : std_logic;
signal \N__20191\ : std_logic;
signal \N__20188\ : std_logic;
signal \N__20185\ : std_logic;
signal \N__20182\ : std_logic;
signal \N__20179\ : std_logic;
signal \N__20178\ : std_logic;
signal \N__20173\ : std_logic;
signal \N__20170\ : std_logic;
signal \N__20169\ : std_logic;
signal \N__20168\ : std_logic;
signal \N__20167\ : std_logic;
signal \N__20166\ : std_logic;
signal \N__20165\ : std_logic;
signal \N__20164\ : std_logic;
signal \N__20161\ : std_logic;
signal \N__20154\ : std_logic;
signal \N__20147\ : std_logic;
signal \N__20144\ : std_logic;
signal \N__20141\ : std_logic;
signal \N__20138\ : std_logic;
signal \N__20135\ : std_logic;
signal \N__20130\ : std_logic;
signal \N__20125\ : std_logic;
signal \N__20122\ : std_logic;
signal \N__20119\ : std_logic;
signal \N__20118\ : std_logic;
signal \N__20115\ : std_logic;
signal \N__20112\ : std_logic;
signal \N__20107\ : std_logic;
signal \N__20106\ : std_logic;
signal \N__20103\ : std_logic;
signal \N__20100\ : std_logic;
signal \N__20095\ : std_logic;
signal \N__20092\ : std_logic;
signal \N__20089\ : std_logic;
signal \N__20086\ : std_logic;
signal \N__20083\ : std_logic;
signal \N__20080\ : std_logic;
signal \N__20077\ : std_logic;
signal \N__20076\ : std_logic;
signal \N__20075\ : std_logic;
signal \N__20074\ : std_logic;
signal \N__20073\ : std_logic;
signal \N__20072\ : std_logic;
signal \N__20071\ : std_logic;
signal \N__20062\ : std_logic;
signal \N__20055\ : std_logic;
signal \N__20052\ : std_logic;
signal \N__20047\ : std_logic;
signal \N__20046\ : std_logic;
signal \N__20045\ : std_logic;
signal \N__20044\ : std_logic;
signal \N__20043\ : std_logic;
signal \N__20042\ : std_logic;
signal \N__20041\ : std_logic;
signal \N__20040\ : std_logic;
signal \N__20031\ : std_logic;
signal \N__20030\ : std_logic;
signal \N__20021\ : std_logic;
signal \N__20018\ : std_logic;
signal \N__20015\ : std_logic;
signal \N__20008\ : std_logic;
signal \N__20007\ : std_logic;
signal \N__20006\ : std_logic;
signal \N__20005\ : std_logic;
signal \N__20002\ : std_logic;
signal \N__19993\ : std_logic;
signal \N__19992\ : std_logic;
signal \N__19991\ : std_logic;
signal \N__19988\ : std_logic;
signal \N__19987\ : std_logic;
signal \N__19984\ : std_logic;
signal \N__19983\ : std_logic;
signal \N__19980\ : std_logic;
signal \N__19979\ : std_logic;
signal \N__19976\ : std_logic;
signal \N__19973\ : std_logic;
signal \N__19966\ : std_logic;
signal \N__19963\ : std_logic;
signal \N__19954\ : std_logic;
signal \N__19951\ : std_logic;
signal \N__19950\ : std_logic;
signal \N__19949\ : std_logic;
signal \N__19948\ : std_logic;
signal \N__19945\ : std_logic;
signal \N__19942\ : std_logic;
signal \N__19939\ : std_logic;
signal \N__19938\ : std_logic;
signal \N__19937\ : std_logic;
signal \N__19934\ : std_logic;
signal \N__19933\ : std_logic;
signal \N__19924\ : std_logic;
signal \N__19923\ : std_logic;
signal \N__19916\ : std_logic;
signal \N__19913\ : std_logic;
signal \N__19910\ : std_logic;
signal \N__19903\ : std_logic;
signal \N__19900\ : std_logic;
signal \N__19897\ : std_logic;
signal \N__19896\ : std_logic;
signal \N__19895\ : std_logic;
signal \N__19894\ : std_logic;
signal \N__19893\ : std_logic;
signal \N__19890\ : std_logic;
signal \N__19889\ : std_logic;
signal \N__19888\ : std_logic;
signal \N__19887\ : std_logic;
signal \N__19886\ : std_logic;
signal \N__19885\ : std_logic;
signal \N__19884\ : std_logic;
signal \N__19883\ : std_logic;
signal \N__19882\ : std_logic;
signal \N__19881\ : std_logic;
signal \N__19880\ : std_logic;
signal \N__19879\ : std_logic;
signal \N__19878\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19876\ : std_logic;
signal \N__19875\ : std_logic;
signal \N__19870\ : std_logic;
signal \N__19865\ : std_logic;
signal \N__19858\ : std_logic;
signal \N__19857\ : std_logic;
signal \N__19856\ : std_logic;
signal \N__19855\ : std_logic;
signal \N__19852\ : std_logic;
signal \N__19851\ : std_logic;
signal \N__19850\ : std_logic;
signal \N__19849\ : std_logic;
signal \N__19848\ : std_logic;
signal \N__19845\ : std_logic;
signal \N__19840\ : std_logic;
signal \N__19835\ : std_logic;
signal \N__19828\ : std_logic;
signal \N__19821\ : std_logic;
signal \N__19820\ : std_logic;
signal \N__19817\ : std_logic;
signal \N__19810\ : std_logic;
signal \N__19807\ : std_logic;
signal \N__19802\ : std_logic;
signal \N__19797\ : std_logic;
signal \N__19790\ : std_logic;
signal \N__19783\ : std_logic;
signal \N__19778\ : std_logic;
signal \N__19773\ : std_logic;
signal \N__19770\ : std_logic;
signal \N__19761\ : std_logic;
signal \N__19758\ : std_logic;
signal \N__19755\ : std_logic;
signal \N__19750\ : std_logic;
signal \N__19741\ : std_logic;
signal \N__19740\ : std_logic;
signal \N__19739\ : std_logic;
signal \N__19738\ : std_logic;
signal \N__19737\ : std_logic;
signal \N__19736\ : std_logic;
signal \N__19733\ : std_logic;
signal \N__19730\ : std_logic;
signal \N__19727\ : std_logic;
signal \N__19726\ : std_logic;
signal \N__19723\ : std_logic;
signal \N__19722\ : std_logic;
signal \N__19713\ : std_logic;
signal \N__19704\ : std_logic;
signal \N__19699\ : std_logic;
signal \N__19696\ : std_logic;
signal \N__19695\ : std_logic;
signal \N__19690\ : std_logic;
signal \N__19687\ : std_logic;
signal \N__19684\ : std_logic;
signal \N__19683\ : std_logic;
signal \N__19682\ : std_logic;
signal \N__19681\ : std_logic;
signal \N__19672\ : std_logic;
signal \N__19671\ : std_logic;
signal \N__19670\ : std_logic;
signal \N__19669\ : std_logic;
signal \N__19668\ : std_logic;
signal \N__19667\ : std_logic;
signal \N__19666\ : std_logic;
signal \N__19665\ : std_logic;
signal \N__19664\ : std_logic;
signal \N__19661\ : std_logic;
signal \N__19660\ : std_logic;
signal \N__19659\ : std_logic;
signal \N__19646\ : std_logic;
signal \N__19645\ : std_logic;
signal \N__19644\ : std_logic;
signal \N__19639\ : std_logic;
signal \N__19636\ : std_logic;
signal \N__19631\ : std_logic;
signal \N__19628\ : std_logic;
signal \N__19623\ : std_logic;
signal \N__19612\ : std_logic;
signal \N__19609\ : std_logic;
signal \N__19608\ : std_logic;
signal \N__19605\ : std_logic;
signal \N__19604\ : std_logic;
signal \N__19603\ : std_logic;
signal \N__19594\ : std_logic;
signal \N__19591\ : std_logic;
signal \N__19590\ : std_logic;
signal \N__19589\ : std_logic;
signal \N__19588\ : std_logic;
signal \N__19587\ : std_logic;
signal \N__19584\ : std_logic;
signal \N__19581\ : std_logic;
signal \N__19576\ : std_logic;
signal \N__19573\ : std_logic;
signal \N__19564\ : std_logic;
signal \N__19563\ : std_logic;
signal \N__19562\ : std_logic;
signal \N__19561\ : std_logic;
signal \N__19560\ : std_logic;
signal \N__19559\ : std_logic;
signal \N__19556\ : std_logic;
signal \N__19549\ : std_logic;
signal \N__19544\ : std_logic;
signal \N__19543\ : std_logic;
signal \N__19536\ : std_logic;
signal \N__19533\ : std_logic;
signal \N__19530\ : std_logic;
signal \N__19527\ : std_logic;
signal \N__19522\ : std_logic;
signal \N__19519\ : std_logic;
signal \N__19516\ : std_logic;
signal \N__19513\ : std_logic;
signal \N__19510\ : std_logic;
signal \N__19507\ : std_logic;
signal \N__19504\ : std_logic;
signal \N__19501\ : std_logic;
signal \N__19498\ : std_logic;
signal \N__19497\ : std_logic;
signal \N__19496\ : std_logic;
signal \N__19495\ : std_logic;
signal \N__19494\ : std_logic;
signal \N__19493\ : std_logic;
signal \N__19492\ : std_logic;
signal \N__19491\ : std_logic;
signal \N__19488\ : std_logic;
signal \N__19487\ : std_logic;
signal \N__19484\ : std_logic;
signal \N__19483\ : std_logic;
signal \N__19480\ : std_logic;
signal \N__19477\ : std_logic;
signal \N__19474\ : std_logic;
signal \N__19473\ : std_logic;
signal \N__19468\ : std_logic;
signal \N__19465\ : std_logic;
signal \N__19460\ : std_logic;
signal \N__19459\ : std_logic;
signal \N__19458\ : std_logic;
signal \N__19453\ : std_logic;
signal \N__19448\ : std_logic;
signal \N__19445\ : std_logic;
signal \N__19442\ : std_logic;
signal \N__19439\ : std_logic;
signal \N__19438\ : std_logic;
signal \N__19437\ : std_logic;
signal \N__19436\ : std_logic;
signal \N__19435\ : std_logic;
signal \N__19432\ : std_logic;
signal \N__19429\ : std_logic;
signal \N__19426\ : std_logic;
signal \N__19425\ : std_logic;
signal \N__19422\ : std_logic;
signal \N__19415\ : std_logic;
signal \N__19410\ : std_logic;
signal \N__19407\ : std_logic;
signal \N__19402\ : std_logic;
signal \N__19399\ : std_logic;
signal \N__19394\ : std_logic;
signal \N__19391\ : std_logic;
signal \N__19386\ : std_logic;
signal \N__19369\ : std_logic;
signal \N__19366\ : std_logic;
signal \N__19363\ : std_logic;
signal \N__19360\ : std_logic;
signal \N__19359\ : std_logic;
signal \N__19358\ : std_logic;
signal \N__19357\ : std_logic;
signal \N__19356\ : std_logic;
signal \N__19355\ : std_logic;
signal \N__19354\ : std_logic;
signal \N__19353\ : std_logic;
signal \N__19344\ : std_logic;
signal \N__19335\ : std_logic;
signal \N__19330\ : std_logic;
signal \N__19327\ : std_logic;
signal \N__19324\ : std_logic;
signal \N__19321\ : std_logic;
signal \N__19318\ : std_logic;
signal \N__19317\ : std_logic;
signal \N__19316\ : std_logic;
signal \N__19315\ : std_logic;
signal \N__19312\ : std_logic;
signal \N__19311\ : std_logic;
signal \N__19310\ : std_logic;
signal \N__19307\ : std_logic;
signal \N__19306\ : std_logic;
signal \N__19305\ : std_logic;
signal \N__19304\ : std_logic;
signal \N__19301\ : std_logic;
signal \N__19298\ : std_logic;
signal \N__19289\ : std_logic;
signal \N__19286\ : std_logic;
signal \N__19277\ : std_logic;
signal \N__19270\ : std_logic;
signal \N__19269\ : std_logic;
signal \N__19268\ : std_logic;
signal \N__19267\ : std_logic;
signal \N__19266\ : std_logic;
signal \N__19265\ : std_logic;
signal \N__19264\ : std_logic;
signal \N__19263\ : std_logic;
signal \N__19254\ : std_logic;
signal \N__19245\ : std_logic;
signal \N__19240\ : std_logic;
signal \N__19239\ : std_logic;
signal \N__19238\ : std_logic;
signal \N__19231\ : std_logic;
signal \N__19228\ : std_logic;
signal \N__19227\ : std_logic;
signal \N__19226\ : std_logic;
signal \N__19219\ : std_logic;
signal \N__19218\ : std_logic;
signal \N__19215\ : std_logic;
signal \N__19212\ : std_logic;
signal \N__19209\ : std_logic;
signal \N__19204\ : std_logic;
signal \N__19201\ : std_logic;
signal \N__19198\ : std_logic;
signal \N__19195\ : std_logic;
signal \N__19192\ : std_logic;
signal \N__19191\ : std_logic;
signal \N__19188\ : std_logic;
signal \N__19187\ : std_logic;
signal \N__19186\ : std_logic;
signal \N__19183\ : std_logic;
signal \N__19176\ : std_logic;
signal \N__19173\ : std_logic;
signal \N__19172\ : std_logic;
signal \N__19171\ : std_logic;
signal \N__19168\ : std_logic;
signal \N__19165\ : std_logic;
signal \N__19162\ : std_logic;
signal \N__19159\ : std_logic;
signal \N__19154\ : std_logic;
signal \N__19147\ : std_logic;
signal \N__19144\ : std_logic;
signal \N__19141\ : std_logic;
signal \N__19140\ : std_logic;
signal \N__19139\ : std_logic;
signal \N__19136\ : std_logic;
signal \N__19131\ : std_logic;
signal \N__19128\ : std_logic;
signal \N__19123\ : std_logic;
signal \N__19120\ : std_logic;
signal \N__19117\ : std_logic;
signal \N__19114\ : std_logic;
signal \N__19111\ : std_logic;
signal \N__19108\ : std_logic;
signal \N__19105\ : std_logic;
signal \N__19102\ : std_logic;
signal \N__19099\ : std_logic;
signal \N__19096\ : std_logic;
signal \N__19093\ : std_logic;
signal \N__19090\ : std_logic;
signal \N__19087\ : std_logic;
signal \N__19084\ : std_logic;
signal \N__19081\ : std_logic;
signal \N__19078\ : std_logic;
signal \N__19075\ : std_logic;
signal \N__19072\ : std_logic;
signal \N__19069\ : std_logic;
signal \N__19068\ : std_logic;
signal \N__19065\ : std_logic;
signal \N__19064\ : std_logic;
signal \N__19063\ : std_logic;
signal \N__19062\ : std_logic;
signal \N__19051\ : std_logic;
signal \N__19050\ : std_logic;
signal \N__19049\ : std_logic;
signal \N__19046\ : std_logic;
signal \N__19041\ : std_logic;
signal \N__19036\ : std_logic;
signal \N__19035\ : std_logic;
signal \N__19034\ : std_logic;
signal \N__19031\ : std_logic;
signal \N__19030\ : std_logic;
signal \N__19027\ : std_logic;
signal \N__19024\ : std_logic;
signal \N__19023\ : std_logic;
signal \N__19018\ : std_logic;
signal \N__19015\ : std_logic;
signal \N__19010\ : std_logic;
signal \N__19007\ : std_logic;
signal \N__19004\ : std_logic;
signal \N__18997\ : std_logic;
signal \N__18994\ : std_logic;
signal \N__18993\ : std_logic;
signal \N__18992\ : std_logic;
signal \N__18991\ : std_logic;
signal \N__18988\ : std_logic;
signal \N__18983\ : std_logic;
signal \N__18980\ : std_logic;
signal \N__18973\ : std_logic;
signal \N__18970\ : std_logic;
signal \N__18969\ : std_logic;
signal \N__18968\ : std_logic;
signal \N__18967\ : std_logic;
signal \N__18964\ : std_logic;
signal \N__18963\ : std_logic;
signal \N__18962\ : std_logic;
signal \N__18955\ : std_logic;
signal \N__18952\ : std_logic;
signal \N__18947\ : std_logic;
signal \N__18940\ : std_logic;
signal \N__18937\ : std_logic;
signal \N__18934\ : std_logic;
signal \N__18933\ : std_logic;
signal \N__18930\ : std_logic;
signal \N__18927\ : std_logic;
signal \N__18924\ : std_logic;
signal \N__18919\ : std_logic;
signal \N__18918\ : std_logic;
signal \N__18915\ : std_logic;
signal \N__18912\ : std_logic;
signal \N__18909\ : std_logic;
signal \N__18906\ : std_logic;
signal \N__18903\ : std_logic;
signal \N__18898\ : std_logic;
signal \N__18895\ : std_logic;
signal \N__18892\ : std_logic;
signal \N__18891\ : std_logic;
signal \N__18888\ : std_logic;
signal \N__18883\ : std_logic;
signal \N__18880\ : std_logic;
signal \N__18879\ : std_logic;
signal \N__18878\ : std_logic;
signal \N__18871\ : std_logic;
signal \N__18868\ : std_logic;
signal \N__18865\ : std_logic;
signal \N__18864\ : std_logic;
signal \N__18863\ : std_logic;
signal \N__18858\ : std_logic;
signal \N__18855\ : std_logic;
signal \N__18852\ : std_logic;
signal \N__18847\ : std_logic;
signal \N__18844\ : std_logic;
signal \N__18841\ : std_logic;
signal \N__18838\ : std_logic;
signal \N__18835\ : std_logic;
signal \N__18832\ : std_logic;
signal \N__18829\ : std_logic;
signal \N__18826\ : std_logic;
signal \N__18823\ : std_logic;
signal \N__18820\ : std_logic;
signal \N__18817\ : std_logic;
signal \N__18814\ : std_logic;
signal \N__18811\ : std_logic;
signal \N__18808\ : std_logic;
signal \N__18805\ : std_logic;
signal \N__18802\ : std_logic;
signal \N__18801\ : std_logic;
signal \N__18800\ : std_logic;
signal \N__18799\ : std_logic;
signal \N__18798\ : std_logic;
signal \N__18787\ : std_logic;
signal \N__18786\ : std_logic;
signal \N__18785\ : std_logic;
signal \N__18782\ : std_logic;
signal \N__18779\ : std_logic;
signal \N__18776\ : std_logic;
signal \N__18775\ : std_logic;
signal \N__18774\ : std_logic;
signal \N__18773\ : std_logic;
signal \N__18772\ : std_logic;
signal \N__18771\ : std_logic;
signal \N__18764\ : std_logic;
signal \N__18761\ : std_logic;
signal \N__18752\ : std_logic;
signal \N__18751\ : std_logic;
signal \N__18750\ : std_logic;
signal \N__18749\ : std_logic;
signal \N__18748\ : std_logic;
signal \N__18745\ : std_logic;
signal \N__18742\ : std_logic;
signal \N__18739\ : std_logic;
signal \N__18734\ : std_logic;
signal \N__18731\ : std_logic;
signal \N__18728\ : std_logic;
signal \N__18715\ : std_logic;
signal \N__18712\ : std_logic;
signal \N__18709\ : std_logic;
signal \N__18706\ : std_logic;
signal \N__18703\ : std_logic;
signal \N__18700\ : std_logic;
signal \N__18697\ : std_logic;
signal \N__18694\ : std_logic;
signal \N__18691\ : std_logic;
signal \N__18690\ : std_logic;
signal \N__18689\ : std_logic;
signal \N__18688\ : std_logic;
signal \N__18685\ : std_logic;
signal \N__18678\ : std_logic;
signal \N__18673\ : std_logic;
signal \N__18672\ : std_logic;
signal \N__18671\ : std_logic;
signal \N__18670\ : std_logic;
signal \N__18667\ : std_logic;
signal \N__18664\ : std_logic;
signal \N__18661\ : std_logic;
signal \N__18656\ : std_logic;
signal \N__18651\ : std_logic;
signal \N__18646\ : std_logic;
signal \N__18645\ : std_logic;
signal \N__18644\ : std_logic;
signal \N__18643\ : std_logic;
signal \N__18640\ : std_logic;
signal \N__18633\ : std_logic;
signal \N__18628\ : std_logic;
signal \N__18625\ : std_logic;
signal \N__18622\ : std_logic;
signal \N__18621\ : std_logic;
signal \N__18620\ : std_logic;
signal \N__18613\ : std_logic;
signal \N__18610\ : std_logic;
signal \N__18609\ : std_logic;
signal \N__18608\ : std_logic;
signal \N__18605\ : std_logic;
signal \N__18604\ : std_logic;
signal \N__18603\ : std_logic;
signal \N__18602\ : std_logic;
signal \N__18601\ : std_logic;
signal \N__18598\ : std_logic;
signal \N__18595\ : std_logic;
signal \N__18594\ : std_logic;
signal \N__18593\ : std_logic;
signal \N__18592\ : std_logic;
signal \N__18585\ : std_logic;
signal \N__18582\ : std_logic;
signal \N__18577\ : std_logic;
signal \N__18568\ : std_logic;
signal \N__18559\ : std_logic;
signal \N__18558\ : std_logic;
signal \N__18557\ : std_logic;
signal \N__18556\ : std_logic;
signal \N__18555\ : std_logic;
signal \N__18554\ : std_logic;
signal \N__18547\ : std_logic;
signal \N__18540\ : std_logic;
signal \N__18535\ : std_logic;
signal \N__18532\ : std_logic;
signal \N__18529\ : std_logic;
signal \N__18526\ : std_logic;
signal \N__18523\ : std_logic;
signal \N__18520\ : std_logic;
signal \N__18517\ : std_logic;
signal \N__18514\ : std_logic;
signal \N__18513\ : std_logic;
signal \N__18508\ : std_logic;
signal \N__18505\ : std_logic;
signal \N__18502\ : std_logic;
signal \N__18501\ : std_logic;
signal \N__18500\ : std_logic;
signal \N__18495\ : std_logic;
signal \N__18492\ : std_logic;
signal \N__18487\ : std_logic;
signal \N__18486\ : std_logic;
signal \N__18483\ : std_logic;
signal \N__18480\ : std_logic;
signal \N__18479\ : std_logic;
signal \N__18476\ : std_logic;
signal \N__18471\ : std_logic;
signal \N__18468\ : std_logic;
signal \N__18463\ : std_logic;
signal \N__18460\ : std_logic;
signal \N__18457\ : std_logic;
signal \N__18454\ : std_logic;
signal \N__18453\ : std_logic;
signal \N__18452\ : std_logic;
signal \N__18451\ : std_logic;
signal \N__18450\ : std_logic;
signal \N__18447\ : std_logic;
signal \N__18440\ : std_logic;
signal \N__18437\ : std_logic;
signal \N__18430\ : std_logic;
signal \N__18429\ : std_logic;
signal \N__18428\ : std_logic;
signal \N__18427\ : std_logic;
signal \N__18424\ : std_logic;
signal \N__18421\ : std_logic;
signal \N__18416\ : std_logic;
signal \N__18409\ : std_logic;
signal \N__18406\ : std_logic;
signal \N__18403\ : std_logic;
signal \N__18400\ : std_logic;
signal \N__18397\ : std_logic;
signal \N__18394\ : std_logic;
signal \N__18391\ : std_logic;
signal \N__18388\ : std_logic;
signal \N__18385\ : std_logic;
signal \N__18382\ : std_logic;
signal \N__18379\ : std_logic;
signal \N__18376\ : std_logic;
signal \N__18375\ : std_logic;
signal \N__18372\ : std_logic;
signal \N__18371\ : std_logic;
signal \N__18368\ : std_logic;
signal \N__18367\ : std_logic;
signal \N__18366\ : std_logic;
signal \N__18361\ : std_logic;
signal \N__18358\ : std_logic;
signal \N__18353\ : std_logic;
signal \N__18348\ : std_logic;
signal \N__18343\ : std_logic;
signal \N__18340\ : std_logic;
signal \N__18337\ : std_logic;
signal \N__18334\ : std_logic;
signal \N__18331\ : std_logic;
signal \N__18328\ : std_logic;
signal \N__18325\ : std_logic;
signal \N__18322\ : std_logic;
signal \N__18321\ : std_logic;
signal \N__18320\ : std_logic;
signal \N__18319\ : std_logic;
signal \N__18318\ : std_logic;
signal \N__18317\ : std_logic;
signal \N__18314\ : std_logic;
signal \N__18311\ : std_logic;
signal \N__18308\ : std_logic;
signal \N__18307\ : std_logic;
signal \N__18306\ : std_logic;
signal \N__18301\ : std_logic;
signal \N__18294\ : std_logic;
signal \N__18287\ : std_logic;
signal \N__18280\ : std_logic;
signal \N__18279\ : std_logic;
signal \N__18278\ : std_logic;
signal \N__18275\ : std_logic;
signal \N__18274\ : std_logic;
signal \N__18273\ : std_logic;
signal \N__18272\ : std_logic;
signal \N__18271\ : std_logic;
signal \N__18270\ : std_logic;
signal \N__18269\ : std_logic;
signal \N__18264\ : std_logic;
signal \N__18261\ : std_logic;
signal \N__18254\ : std_logic;
signal \N__18247\ : std_logic;
signal \N__18238\ : std_logic;
signal \N__18237\ : std_logic;
signal \N__18236\ : std_logic;
signal \N__18235\ : std_logic;
signal \N__18234\ : std_logic;
signal \N__18233\ : std_logic;
signal \N__18232\ : std_logic;
signal \N__18227\ : std_logic;
signal \N__18226\ : std_logic;
signal \N__18225\ : std_logic;
signal \N__18224\ : std_logic;
signal \N__18217\ : std_logic;
signal \N__18212\ : std_logic;
signal \N__18209\ : std_logic;
signal \N__18204\ : std_logic;
signal \N__18201\ : std_logic;
signal \N__18190\ : std_logic;
signal \N__18187\ : std_logic;
signal \N__18186\ : std_logic;
signal \N__18183\ : std_logic;
signal \N__18180\ : std_logic;
signal \N__18179\ : std_logic;
signal \N__18176\ : std_logic;
signal \N__18175\ : std_logic;
signal \N__18174\ : std_logic;
signal \N__18173\ : std_logic;
signal \N__18172\ : std_logic;
signal \N__18171\ : std_logic;
signal \N__18168\ : std_logic;
signal \N__18165\ : std_logic;
signal \N__18162\ : std_logic;
signal \N__18155\ : std_logic;
signal \N__18152\ : std_logic;
signal \N__18149\ : std_logic;
signal \N__18146\ : std_logic;
signal \N__18143\ : std_logic;
signal \N__18130\ : std_logic;
signal \N__18127\ : std_logic;
signal \N__18124\ : std_logic;
signal \N__18121\ : std_logic;
signal \N__18118\ : std_logic;
signal \N__18115\ : std_logic;
signal \N__18112\ : std_logic;
signal \N__18111\ : std_logic;
signal \N__18108\ : std_logic;
signal \N__18105\ : std_logic;
signal \N__18102\ : std_logic;
signal \N__18099\ : std_logic;
signal \N__18096\ : std_logic;
signal \N__18093\ : std_logic;
signal \N__18088\ : std_logic;
signal \N__18085\ : std_logic;
signal \N__18084\ : std_logic;
signal \N__18081\ : std_logic;
signal \N__18078\ : std_logic;
signal \N__18075\ : std_logic;
signal \N__18070\ : std_logic;
signal \N__18067\ : std_logic;
signal \N__18064\ : std_logic;
signal \N__18063\ : std_logic;
signal \N__18062\ : std_logic;
signal \N__18061\ : std_logic;
signal \N__18060\ : std_logic;
signal \N__18059\ : std_logic;
signal \N__18058\ : std_logic;
signal \N__18057\ : std_logic;
signal \N__18056\ : std_logic;
signal \N__18055\ : std_logic;
signal \N__18054\ : std_logic;
signal \N__18053\ : std_logic;
signal \N__18048\ : std_logic;
signal \N__18047\ : std_logic;
signal \N__18046\ : std_logic;
signal \N__18043\ : std_logic;
signal \N__18042\ : std_logic;
signal \N__18041\ : std_logic;
signal \N__18038\ : std_logic;
signal \N__18031\ : std_logic;
signal \N__18026\ : std_logic;
signal \N__18023\ : std_logic;
signal \N__18018\ : std_logic;
signal \N__18015\ : std_logic;
signal \N__18014\ : std_logic;
signal \N__18013\ : std_logic;
signal \N__18010\ : std_logic;
signal \N__18009\ : std_logic;
signal \N__18008\ : std_logic;
signal \N__18007\ : std_logic;
signal \N__18006\ : std_logic;
signal \N__18003\ : std_logic;
signal \N__18000\ : std_logic;
signal \N__17997\ : std_logic;
signal \N__17994\ : std_logic;
signal \N__17987\ : std_logic;
signal \N__17982\ : std_logic;
signal \N__17979\ : std_logic;
signal \N__17976\ : std_logic;
signal \N__17973\ : std_logic;
signal \N__17966\ : std_logic;
signal \N__17963\ : std_logic;
signal \N__17960\ : std_logic;
signal \N__17951\ : std_logic;
signal \N__17946\ : std_logic;
signal \N__17929\ : std_logic;
signal \N__17928\ : std_logic;
signal \N__17927\ : std_logic;
signal \N__17926\ : std_logic;
signal \N__17925\ : std_logic;
signal \N__17924\ : std_logic;
signal \N__17921\ : std_logic;
signal \N__17920\ : std_logic;
signal \N__17919\ : std_logic;
signal \N__17918\ : std_logic;
signal \N__17917\ : std_logic;
signal \N__17916\ : std_logic;
signal \N__17915\ : std_logic;
signal \N__17914\ : std_logic;
signal \N__17913\ : std_logic;
signal \N__17912\ : std_logic;
signal \N__17911\ : std_logic;
signal \N__17910\ : std_logic;
signal \N__17907\ : std_logic;
signal \N__17906\ : std_logic;
signal \N__17905\ : std_logic;
signal \N__17904\ : std_logic;
signal \N__17895\ : std_logic;
signal \N__17894\ : std_logic;
signal \N__17893\ : std_logic;
signal \N__17892\ : std_logic;
signal \N__17889\ : std_logic;
signal \N__17888\ : std_logic;
signal \N__17887\ : std_logic;
signal \N__17886\ : std_logic;
signal \N__17883\ : std_logic;
signal \N__17876\ : std_logic;
signal \N__17873\ : std_logic;
signal \N__17870\ : std_logic;
signal \N__17863\ : std_logic;
signal \N__17862\ : std_logic;
signal \N__17861\ : std_logic;
signal \N__17860\ : std_logic;
signal \N__17859\ : std_logic;
signal \N__17856\ : std_logic;
signal \N__17855\ : std_logic;
signal \N__17854\ : std_logic;
signal \N__17851\ : std_logic;
signal \N__17848\ : std_logic;
signal \N__17841\ : std_logic;
signal \N__17838\ : std_logic;
signal \N__17835\ : std_logic;
signal \N__17832\ : std_logic;
signal \N__17829\ : std_logic;
signal \N__17828\ : std_logic;
signal \N__17825\ : std_logic;
signal \N__17818\ : std_logic;
signal \N__17811\ : std_logic;
signal \N__17806\ : std_logic;
signal \N__17803\ : std_logic;
signal \N__17800\ : std_logic;
signal \N__17795\ : std_logic;
signal \N__17792\ : std_logic;
signal \N__17785\ : std_logic;
signal \N__17778\ : std_logic;
signal \N__17773\ : std_logic;
signal \N__17770\ : std_logic;
signal \N__17767\ : std_logic;
signal \N__17760\ : std_logic;
signal \N__17753\ : std_logic;
signal \N__17750\ : std_logic;
signal \N__17745\ : std_logic;
signal \N__17742\ : std_logic;
signal \N__17725\ : std_logic;
signal \N__17724\ : std_logic;
signal \N__17721\ : std_logic;
signal \N__17718\ : std_logic;
signal \N__17713\ : std_logic;
signal \N__17710\ : std_logic;
signal \N__17707\ : std_logic;
signal \N__17704\ : std_logic;
signal \N__17701\ : std_logic;
signal \N__17698\ : std_logic;
signal \N__17697\ : std_logic;
signal \N__17696\ : std_logic;
signal \N__17695\ : std_logic;
signal \N__17694\ : std_logic;
signal \N__17691\ : std_logic;
signal \N__17688\ : std_logic;
signal \N__17683\ : std_logic;
signal \N__17680\ : std_logic;
signal \N__17671\ : std_logic;
signal \N__17668\ : std_logic;
signal \N__17667\ : std_logic;
signal \N__17664\ : std_logic;
signal \N__17661\ : std_logic;
signal \N__17660\ : std_logic;
signal \N__17657\ : std_logic;
signal \N__17654\ : std_logic;
signal \N__17651\ : std_logic;
signal \N__17650\ : std_logic;
signal \N__17649\ : std_logic;
signal \N__17642\ : std_logic;
signal \N__17639\ : std_logic;
signal \N__17636\ : std_logic;
signal \N__17629\ : std_logic;
signal \N__17626\ : std_logic;
signal \N__17623\ : std_logic;
signal \N__17620\ : std_logic;
signal \N__17617\ : std_logic;
signal \N__17616\ : std_logic;
signal \N__17613\ : std_logic;
signal \N__17610\ : std_logic;
signal \N__17607\ : std_logic;
signal \N__17602\ : std_logic;
signal \N__17599\ : std_logic;
signal \N__17596\ : std_logic;
signal \N__17593\ : std_logic;
signal \N__17590\ : std_logic;
signal \N__17587\ : std_logic;
signal \N__17584\ : std_logic;
signal \N__17581\ : std_logic;
signal \N__17578\ : std_logic;
signal \N__17575\ : std_logic;
signal \N__17572\ : std_logic;
signal \N__17571\ : std_logic;
signal \N__17568\ : std_logic;
signal \N__17567\ : std_logic;
signal \N__17566\ : std_logic;
signal \N__17565\ : std_logic;
signal \N__17562\ : std_logic;
signal \N__17559\ : std_logic;
signal \N__17554\ : std_logic;
signal \N__17553\ : std_logic;
signal \N__17552\ : std_logic;
signal \N__17549\ : std_logic;
signal \N__17548\ : std_logic;
signal \N__17547\ : std_logic;
signal \N__17546\ : std_logic;
signal \N__17543\ : std_logic;
signal \N__17538\ : std_logic;
signal \N__17533\ : std_logic;
signal \N__17532\ : std_logic;
signal \N__17527\ : std_logic;
signal \N__17526\ : std_logic;
signal \N__17521\ : std_logic;
signal \N__17516\ : std_logic;
signal \N__17513\ : std_logic;
signal \N__17510\ : std_logic;
signal \N__17507\ : std_logic;
signal \N__17504\ : std_logic;
signal \N__17491\ : std_logic;
signal \N__17488\ : std_logic;
signal \N__17485\ : std_logic;
signal \N__17482\ : std_logic;
signal \N__17479\ : std_logic;
signal \N__17476\ : std_logic;
signal \N__17473\ : std_logic;
signal \N__17472\ : std_logic;
signal \N__17469\ : std_logic;
signal \N__17466\ : std_logic;
signal \N__17461\ : std_logic;
signal \N__17458\ : std_logic;
signal \N__17455\ : std_logic;
signal \N__17452\ : std_logic;
signal \N__17449\ : std_logic;
signal \N__17446\ : std_logic;
signal \N__17443\ : std_logic;
signal \N__17442\ : std_logic;
signal \N__17437\ : std_logic;
signal \N__17434\ : std_logic;
signal \N__17431\ : std_logic;
signal \N__17428\ : std_logic;
signal \N__17425\ : std_logic;
signal \N__17422\ : std_logic;
signal \N__17419\ : std_logic;
signal \N__17416\ : std_logic;
signal \N__17415\ : std_logic;
signal \N__17412\ : std_logic;
signal \N__17409\ : std_logic;
signal \N__17404\ : std_logic;
signal \N__17401\ : std_logic;
signal \N__17398\ : std_logic;
signal \N__17395\ : std_logic;
signal \N__17394\ : std_logic;
signal \N__17391\ : std_logic;
signal \N__17388\ : std_logic;
signal \N__17383\ : std_logic;
signal \N__17380\ : std_logic;
signal \N__17377\ : std_logic;
signal \N__17374\ : std_logic;
signal \N__17371\ : std_logic;
signal \N__17368\ : std_logic;
signal \N__17365\ : std_logic;
signal \N__17364\ : std_logic;
signal \N__17359\ : std_logic;
signal \N__17356\ : std_logic;
signal \N__17355\ : std_logic;
signal \N__17352\ : std_logic;
signal \N__17351\ : std_logic;
signal \N__17350\ : std_logic;
signal \N__17345\ : std_logic;
signal \N__17340\ : std_logic;
signal \N__17335\ : std_logic;
signal \N__17332\ : std_logic;
signal \N__17331\ : std_logic;
signal \N__17328\ : std_logic;
signal \N__17325\ : std_logic;
signal \N__17322\ : std_logic;
signal \N__17319\ : std_logic;
signal \N__17316\ : std_logic;
signal \N__17313\ : std_logic;
signal \N__17308\ : std_logic;
signal \N__17307\ : std_logic;
signal \N__17306\ : std_logic;
signal \N__17305\ : std_logic;
signal \N__17304\ : std_logic;
signal \N__17303\ : std_logic;
signal \N__17302\ : std_logic;
signal \N__17293\ : std_logic;
signal \N__17290\ : std_logic;
signal \N__17285\ : std_logic;
signal \N__17282\ : std_logic;
signal \N__17277\ : std_logic;
signal \N__17274\ : std_logic;
signal \N__17271\ : std_logic;
signal \N__17266\ : std_logic;
signal \N__17265\ : std_logic;
signal \N__17264\ : std_logic;
signal \N__17263\ : std_logic;
signal \N__17262\ : std_logic;
signal \N__17261\ : std_logic;
signal \N__17260\ : std_logic;
signal \N__17259\ : std_logic;
signal \N__17258\ : std_logic;
signal \N__17257\ : std_logic;
signal \N__17254\ : std_logic;
signal \N__17247\ : std_logic;
signal \N__17244\ : std_logic;
signal \N__17241\ : std_logic;
signal \N__17232\ : std_logic;
signal \N__17231\ : std_logic;
signal \N__17230\ : std_logic;
signal \N__17225\ : std_logic;
signal \N__17222\ : std_logic;
signal \N__17221\ : std_logic;
signal \N__17216\ : std_logic;
signal \N__17213\ : std_logic;
signal \N__17210\ : std_logic;
signal \N__17205\ : std_logic;
signal \N__17202\ : std_logic;
signal \N__17199\ : std_logic;
signal \N__17194\ : std_logic;
signal \N__17185\ : std_logic;
signal \N__17184\ : std_logic;
signal \N__17183\ : std_logic;
signal \N__17182\ : std_logic;
signal \N__17181\ : std_logic;
signal \N__17178\ : std_logic;
signal \N__17175\ : std_logic;
signal \N__17172\ : std_logic;
signal \N__17169\ : std_logic;
signal \N__17166\ : std_logic;
signal \N__17161\ : std_logic;
signal \N__17156\ : std_logic;
signal \N__17153\ : std_logic;
signal \N__17148\ : std_logic;
signal \N__17145\ : std_logic;
signal \N__17142\ : std_logic;
signal \N__17137\ : std_logic;
signal \N__17134\ : std_logic;
signal \N__17131\ : std_logic;
signal \N__17128\ : std_logic;
signal \N__17125\ : std_logic;
signal \N__17122\ : std_logic;
signal \N__17119\ : std_logic;
signal \N__17116\ : std_logic;
signal \N__17113\ : std_logic;
signal \N__17112\ : std_logic;
signal \N__17109\ : std_logic;
signal \N__17106\ : std_logic;
signal \N__17103\ : std_logic;
signal \N__17100\ : std_logic;
signal \N__17099\ : std_logic;
signal \N__17094\ : std_logic;
signal \N__17091\ : std_logic;
signal \N__17088\ : std_logic;
signal \N__17083\ : std_logic;
signal \N__17080\ : std_logic;
signal \N__17077\ : std_logic;
signal \N__17074\ : std_logic;
signal \N__17071\ : std_logic;
signal \N__17068\ : std_logic;
signal \N__17065\ : std_logic;
signal \N__17062\ : std_logic;
signal \N__17059\ : std_logic;
signal \N__17056\ : std_logic;
signal \N__17053\ : std_logic;
signal \N__17050\ : std_logic;
signal \N__17047\ : std_logic;
signal \N__17044\ : std_logic;
signal \N__17043\ : std_logic;
signal \N__17042\ : std_logic;
signal \N__17041\ : std_logic;
signal \N__17040\ : std_logic;
signal \N__17039\ : std_logic;
signal \N__17038\ : std_logic;
signal \N__17037\ : std_logic;
signal \N__17034\ : std_logic;
signal \N__17033\ : std_logic;
signal \N__17032\ : std_logic;
signal \N__17023\ : std_logic;
signal \N__17012\ : std_logic;
signal \N__17009\ : std_logic;
signal \N__17002\ : std_logic;
signal \N__17001\ : std_logic;
signal \N__17000\ : std_logic;
signal \N__16999\ : std_logic;
signal \N__16998\ : std_logic;
signal \N__16995\ : std_logic;
signal \N__16994\ : std_logic;
signal \N__16991\ : std_logic;
signal \N__16988\ : std_logic;
signal \N__16987\ : std_logic;
signal \N__16984\ : std_logic;
signal \N__16983\ : std_logic;
signal \N__16980\ : std_logic;
signal \N__16979\ : std_logic;
signal \N__16970\ : std_logic;
signal \N__16967\ : std_logic;
signal \N__16958\ : std_logic;
signal \N__16951\ : std_logic;
signal \N__16948\ : std_logic;
signal \N__16945\ : std_logic;
signal \N__16942\ : std_logic;
signal \N__16941\ : std_logic;
signal \N__16940\ : std_logic;
signal \N__16939\ : std_logic;
signal \N__16938\ : std_logic;
signal \N__16937\ : std_logic;
signal \N__16936\ : std_logic;
signal \N__16935\ : std_logic;
signal \N__16934\ : std_logic;
signal \N__16925\ : std_logic;
signal \N__16922\ : std_logic;
signal \N__16913\ : std_logic;
signal \N__16906\ : std_logic;
signal \N__16903\ : std_logic;
signal \N__16900\ : std_logic;
signal \N__16897\ : std_logic;
signal \N__16894\ : std_logic;
signal \N__16891\ : std_logic;
signal \N__16888\ : std_logic;
signal \N__16885\ : std_logic;
signal \N__16882\ : std_logic;
signal \N__16879\ : std_logic;
signal \N__16876\ : std_logic;
signal \N__16873\ : std_logic;
signal \N__16870\ : std_logic;
signal \N__16867\ : std_logic;
signal \N__16864\ : std_logic;
signal \N__16861\ : std_logic;
signal \N__16858\ : std_logic;
signal \N__16857\ : std_logic;
signal \N__16852\ : std_logic;
signal \N__16849\ : std_logic;
signal \N__16846\ : std_logic;
signal \N__16843\ : std_logic;
signal \N__16840\ : std_logic;
signal \N__16837\ : std_logic;
signal \N__16834\ : std_logic;
signal \N__16833\ : std_logic;
signal \N__16828\ : std_logic;
signal \N__16825\ : std_logic;
signal \N__16822\ : std_logic;
signal \N__16819\ : std_logic;
signal \N__16816\ : std_logic;
signal \N__16813\ : std_logic;
signal \N__16810\ : std_logic;
signal \N__16807\ : std_logic;
signal \N__16804\ : std_logic;
signal \N__16801\ : std_logic;
signal \N__16798\ : std_logic;
signal \N__16795\ : std_logic;
signal \N__16792\ : std_logic;
signal \N__16789\ : std_logic;
signal \N__16788\ : std_logic;
signal \N__16787\ : std_logic;
signal \N__16786\ : std_logic;
signal \N__16781\ : std_logic;
signal \N__16780\ : std_logic;
signal \N__16779\ : std_logic;
signal \N__16778\ : std_logic;
signal \N__16777\ : std_logic;
signal \N__16772\ : std_logic;
signal \N__16771\ : std_logic;
signal \N__16770\ : std_logic;
signal \N__16769\ : std_logic;
signal \N__16768\ : std_logic;
signal \N__16767\ : std_logic;
signal \N__16764\ : std_logic;
signal \N__16761\ : std_logic;
signal \N__16758\ : std_logic;
signal \N__16757\ : std_logic;
signal \N__16756\ : std_logic;
signal \N__16751\ : std_logic;
signal \N__16748\ : std_logic;
signal \N__16745\ : std_logic;
signal \N__16740\ : std_logic;
signal \N__16737\ : std_logic;
signal \N__16734\ : std_logic;
signal \N__16731\ : std_logic;
signal \N__16728\ : std_logic;
signal \N__16721\ : std_logic;
signal \N__16702\ : std_logic;
signal \N__16699\ : std_logic;
signal \N__16696\ : std_logic;
signal \N__16693\ : std_logic;
signal \N__16690\ : std_logic;
signal \N__16687\ : std_logic;
signal \N__16684\ : std_logic;
signal \N__16681\ : std_logic;
signal \N__16678\ : std_logic;
signal \N__16675\ : std_logic;
signal \N__16672\ : std_logic;
signal \N__16669\ : std_logic;
signal \N__16666\ : std_logic;
signal \N__16663\ : std_logic;
signal \N__16660\ : std_logic;
signal \N__16657\ : std_logic;
signal \N__16654\ : std_logic;
signal \N__16651\ : std_logic;
signal \N__16648\ : std_logic;
signal \N__16645\ : std_logic;
signal \N__16644\ : std_logic;
signal \N__16643\ : std_logic;
signal \N__16642\ : std_logic;
signal \N__16641\ : std_logic;
signal \N__16640\ : std_logic;
signal \N__16639\ : std_logic;
signal \N__16636\ : std_logic;
signal \N__16633\ : std_logic;
signal \N__16628\ : std_logic;
signal \N__16627\ : std_logic;
signal \N__16622\ : std_logic;
signal \N__16619\ : std_logic;
signal \N__16618\ : std_logic;
signal \N__16617\ : std_logic;
signal \N__16616\ : std_logic;
signal \N__16613\ : std_logic;
signal \N__16608\ : std_logic;
signal \N__16605\ : std_logic;
signal \N__16604\ : std_logic;
signal \N__16601\ : std_logic;
signal \N__16598\ : std_logic;
signal \N__16595\ : std_logic;
signal \N__16590\ : std_logic;
signal \N__16583\ : std_logic;
signal \N__16580\ : std_logic;
signal \N__16577\ : std_logic;
signal \N__16564\ : std_logic;
signal \N__16561\ : std_logic;
signal \N__16558\ : std_logic;
signal \N__16555\ : std_logic;
signal \N__16552\ : std_logic;
signal \N__16549\ : std_logic;
signal \N__16546\ : std_logic;
signal \N__16545\ : std_logic;
signal \N__16544\ : std_logic;
signal \N__16543\ : std_logic;
signal \N__16540\ : std_logic;
signal \N__16537\ : std_logic;
signal \N__16534\ : std_logic;
signal \N__16533\ : std_logic;
signal \N__16530\ : std_logic;
signal \N__16525\ : std_logic;
signal \N__16520\ : std_logic;
signal \N__16513\ : std_logic;
signal \N__16512\ : std_logic;
signal \N__16507\ : std_logic;
signal \N__16506\ : std_logic;
signal \N__16505\ : std_logic;
signal \N__16504\ : std_logic;
signal \N__16501\ : std_logic;
signal \N__16500\ : std_logic;
signal \N__16499\ : std_logic;
signal \N__16498\ : std_logic;
signal \N__16495\ : std_logic;
signal \N__16492\ : std_logic;
signal \N__16489\ : std_logic;
signal \N__16486\ : std_logic;
signal \N__16481\ : std_logic;
signal \N__16478\ : std_logic;
signal \N__16465\ : std_logic;
signal \N__16462\ : std_logic;
signal \N__16461\ : std_logic;
signal \N__16458\ : std_logic;
signal \N__16455\ : std_logic;
signal \N__16452\ : std_logic;
signal \N__16447\ : std_logic;
signal \N__16446\ : std_logic;
signal \N__16443\ : std_logic;
signal \N__16442\ : std_logic;
signal \N__16441\ : std_logic;
signal \N__16440\ : std_logic;
signal \N__16437\ : std_logic;
signal \N__16434\ : std_logic;
signal \N__16433\ : std_logic;
signal \N__16430\ : std_logic;
signal \N__16425\ : std_logic;
signal \N__16422\ : std_logic;
signal \N__16419\ : std_logic;
signal \N__16416\ : std_logic;
signal \N__16413\ : std_logic;
signal \N__16402\ : std_logic;
signal \N__16399\ : std_logic;
signal \N__16398\ : std_logic;
signal \N__16397\ : std_logic;
signal \N__16392\ : std_logic;
signal \N__16389\ : std_logic;
signal \N__16388\ : std_logic;
signal \N__16385\ : std_logic;
signal \N__16380\ : std_logic;
signal \N__16375\ : std_logic;
signal \N__16374\ : std_logic;
signal \N__16371\ : std_logic;
signal \N__16368\ : std_logic;
signal \N__16365\ : std_logic;
signal \N__16364\ : std_logic;
signal \N__16363\ : std_logic;
signal \N__16362\ : std_logic;
signal \N__16361\ : std_logic;
signal \N__16358\ : std_logic;
signal \N__16355\ : std_logic;
signal \N__16346\ : std_logic;
signal \N__16339\ : std_logic;
signal \N__16336\ : std_logic;
signal \N__16333\ : std_logic;
signal \N__16332\ : std_logic;
signal \N__16331\ : std_logic;
signal \N__16330\ : std_logic;
signal \N__16329\ : std_logic;
signal \N__16326\ : std_logic;
signal \N__16323\ : std_logic;
signal \N__16316\ : std_logic;
signal \N__16311\ : std_logic;
signal \N__16306\ : std_logic;
signal \N__16303\ : std_logic;
signal \N__16300\ : std_logic;
signal \N__16297\ : std_logic;
signal \N__16294\ : std_logic;
signal \N__16291\ : std_logic;
signal \N__16288\ : std_logic;
signal \N__16285\ : std_logic;
signal \N__16282\ : std_logic;
signal \N__16279\ : std_logic;
signal \N__16276\ : std_logic;
signal \N__16275\ : std_logic;
signal \N__16274\ : std_logic;
signal \N__16273\ : std_logic;
signal \N__16272\ : std_logic;
signal \N__16271\ : std_logic;
signal \N__16268\ : std_logic;
signal \N__16267\ : std_logic;
signal \N__16260\ : std_logic;
signal \N__16259\ : std_logic;
signal \N__16258\ : std_logic;
signal \N__16257\ : std_logic;
signal \N__16256\ : std_logic;
signal \N__16255\ : std_logic;
signal \N__16254\ : std_logic;
signal \N__16253\ : std_logic;
signal \N__16252\ : std_logic;
signal \N__16251\ : std_logic;
signal \N__16250\ : std_logic;
signal \N__16247\ : std_logic;
signal \N__16244\ : std_logic;
signal \N__16241\ : std_logic;
signal \N__16238\ : std_logic;
signal \N__16235\ : std_logic;
signal \N__16232\ : std_logic;
signal \N__16227\ : std_logic;
signal \N__16218\ : std_logic;
signal \N__16209\ : std_logic;
signal \N__16192\ : std_logic;
signal \N__16189\ : std_logic;
signal \N__16186\ : std_logic;
signal \N__16183\ : std_logic;
signal \N__16180\ : std_logic;
signal \N__16177\ : std_logic;
signal \N__16174\ : std_logic;
signal \N__16173\ : std_logic;
signal \N__16172\ : std_logic;
signal \N__16169\ : std_logic;
signal \N__16164\ : std_logic;
signal \N__16159\ : std_logic;
signal \N__16156\ : std_logic;
signal \N__16155\ : std_logic;
signal \N__16152\ : std_logic;
signal \N__16151\ : std_logic;
signal \N__16150\ : std_logic;
signal \N__16147\ : std_logic;
signal \N__16144\ : std_logic;
signal \N__16137\ : std_logic;
signal \N__16132\ : std_logic;
signal \N__16131\ : std_logic;
signal \N__16130\ : std_logic;
signal \N__16129\ : std_logic;
signal \N__16122\ : std_logic;
signal \N__16121\ : std_logic;
signal \N__16120\ : std_logic;
signal \N__16119\ : std_logic;
signal \N__16118\ : std_logic;
signal \N__16115\ : std_logic;
signal \N__16112\ : std_logic;
signal \N__16111\ : std_logic;
signal \N__16110\ : std_logic;
signal \N__16109\ : std_logic;
signal \N__16108\ : std_logic;
signal \N__16105\ : std_logic;
signal \N__16104\ : std_logic;
signal \N__16103\ : std_logic;
signal \N__16098\ : std_logic;
signal \N__16095\ : std_logic;
signal \N__16092\ : std_logic;
signal \N__16089\ : std_logic;
signal \N__16084\ : std_logic;
signal \N__16081\ : std_logic;
signal \N__16072\ : std_logic;
signal \N__16057\ : std_logic;
signal \N__16054\ : std_logic;
signal \N__16053\ : std_logic;
signal \N__16052\ : std_logic;
signal \N__16047\ : std_logic;
signal \N__16044\ : std_logic;
signal \N__16041\ : std_logic;
signal \N__16038\ : std_logic;
signal \N__16033\ : std_logic;
signal \N__16030\ : std_logic;
signal \N__16029\ : std_logic;
signal \N__16026\ : std_logic;
signal \N__16023\ : std_logic;
signal \N__16020\ : std_logic;
signal \N__16015\ : std_logic;
signal \N__16012\ : std_logic;
signal \N__16009\ : std_logic;
signal \N__16006\ : std_logic;
signal \N__16005\ : std_logic;
signal \N__16004\ : std_logic;
signal \N__16001\ : std_logic;
signal \N__15996\ : std_logic;
signal \N__15993\ : std_logic;
signal \N__15988\ : std_logic;
signal \N__15985\ : std_logic;
signal \N__15982\ : std_logic;
signal \N__15979\ : std_logic;
signal \N__15978\ : std_logic;
signal \N__15977\ : std_logic;
signal \N__15976\ : std_logic;
signal \N__15975\ : std_logic;
signal \N__15974\ : std_logic;
signal \N__15973\ : std_logic;
signal \N__15972\ : std_logic;
signal \N__15955\ : std_logic;
signal \N__15954\ : std_logic;
signal \N__15951\ : std_logic;
signal \N__15948\ : std_logic;
signal \N__15943\ : std_logic;
signal \N__15942\ : std_logic;
signal \N__15941\ : std_logic;
signal \N__15938\ : std_logic;
signal \N__15935\ : std_logic;
signal \N__15932\ : std_logic;
signal \N__15931\ : std_logic;
signal \N__15930\ : std_logic;
signal \N__15929\ : std_logic;
signal \N__15928\ : std_logic;
signal \N__15927\ : std_logic;
signal \N__15926\ : std_logic;
signal \N__15925\ : std_logic;
signal \N__15924\ : std_logic;
signal \N__15923\ : std_logic;
signal \N__15922\ : std_logic;
signal \N__15921\ : std_logic;
signal \N__15920\ : std_logic;
signal \N__15919\ : std_logic;
signal \N__15902\ : std_logic;
signal \N__15897\ : std_logic;
signal \N__15892\ : std_logic;
signal \N__15887\ : std_logic;
signal \N__15882\ : std_logic;
signal \N__15871\ : std_logic;
signal \N__15870\ : std_logic;
signal \N__15867\ : std_logic;
signal \N__15864\ : std_logic;
signal \N__15861\ : std_logic;
signal \N__15858\ : std_logic;
signal \N__15855\ : std_logic;
signal \N__15852\ : std_logic;
signal \N__15849\ : std_logic;
signal \N__15844\ : std_logic;
signal \N__15843\ : std_logic;
signal \N__15842\ : std_logic;
signal \N__15839\ : std_logic;
signal \N__15838\ : std_logic;
signal \N__15837\ : std_logic;
signal \N__15836\ : std_logic;
signal \N__15835\ : std_logic;
signal \N__15832\ : std_logic;
signal \N__15829\ : std_logic;
signal \N__15826\ : std_logic;
signal \N__15817\ : std_logic;
signal \N__15814\ : std_logic;
signal \N__15805\ : std_logic;
signal \N__15804\ : std_logic;
signal \N__15803\ : std_logic;
signal \N__15800\ : std_logic;
signal \N__15797\ : std_logic;
signal \N__15796\ : std_logic;
signal \N__15795\ : std_logic;
signal \N__15794\ : std_logic;
signal \N__15793\ : std_logic;
signal \N__15790\ : std_logic;
signal \N__15787\ : std_logic;
signal \N__15784\ : std_logic;
signal \N__15781\ : std_logic;
signal \N__15778\ : std_logic;
signal \N__15773\ : std_logic;
signal \N__15760\ : std_logic;
signal \N__15757\ : std_logic;
signal \N__15754\ : std_logic;
signal \N__15751\ : std_logic;
signal \N__15748\ : std_logic;
signal \N__15745\ : std_logic;
signal \N__15744\ : std_logic;
signal \N__15741\ : std_logic;
signal \N__15740\ : std_logic;
signal \N__15737\ : std_logic;
signal \N__15730\ : std_logic;
signal \N__15727\ : std_logic;
signal \N__15724\ : std_logic;
signal \N__15721\ : std_logic;
signal \N__15720\ : std_logic;
signal \N__15717\ : std_logic;
signal \N__15712\ : std_logic;
signal \N__15709\ : std_logic;
signal \N__15706\ : std_logic;
signal \N__15703\ : std_logic;
signal \N__15700\ : std_logic;
signal \N__15699\ : std_logic;
signal \N__15696\ : std_logic;
signal \N__15691\ : std_logic;
signal \N__15688\ : std_logic;
signal \N__15685\ : std_logic;
signal \N__15682\ : std_logic;
signal \N__15681\ : std_logic;
signal \N__15676\ : std_logic;
signal \N__15673\ : std_logic;
signal \N__15670\ : std_logic;
signal \N__15669\ : std_logic;
signal \N__15666\ : std_logic;
signal \N__15663\ : std_logic;
signal \N__15658\ : std_logic;
signal \N__15655\ : std_logic;
signal \N__15652\ : std_logic;
signal \N__15649\ : std_logic;
signal \N__15646\ : std_logic;
signal \N__15643\ : std_logic;
signal \N__15640\ : std_logic;
signal \N__15637\ : std_logic;
signal \N__15636\ : std_logic;
signal \N__15633\ : std_logic;
signal \N__15630\ : std_logic;
signal \N__15625\ : std_logic;
signal \N__15624\ : std_logic;
signal \N__15621\ : std_logic;
signal \N__15620\ : std_logic;
signal \N__15619\ : std_logic;
signal \N__15616\ : std_logic;
signal \N__15613\ : std_logic;
signal \N__15608\ : std_logic;
signal \N__15601\ : std_logic;
signal \N__15598\ : std_logic;
signal \N__15595\ : std_logic;
signal \N__15592\ : std_logic;
signal \N__15589\ : std_logic;
signal \N__15586\ : std_logic;
signal \N__15583\ : std_logic;
signal \N__15582\ : std_logic;
signal \N__15579\ : std_logic;
signal \N__15576\ : std_logic;
signal \N__15575\ : std_logic;
signal \N__15572\ : std_logic;
signal \N__15569\ : std_logic;
signal \N__15568\ : std_logic;
signal \N__15565\ : std_logic;
signal \N__15562\ : std_logic;
signal \N__15559\ : std_logic;
signal \N__15554\ : std_logic;
signal \N__15551\ : std_logic;
signal \N__15544\ : std_logic;
signal \N__15541\ : std_logic;
signal \N__15538\ : std_logic;
signal \N__15537\ : std_logic;
signal \N__15534\ : std_logic;
signal \N__15531\ : std_logic;
signal \N__15528\ : std_logic;
signal \N__15525\ : std_logic;
signal \N__15522\ : std_logic;
signal \N__15517\ : std_logic;
signal \N__15514\ : std_logic;
signal \N__15513\ : std_logic;
signal \N__15510\ : std_logic;
signal \N__15507\ : std_logic;
signal \N__15504\ : std_logic;
signal \N__15501\ : std_logic;
signal \N__15496\ : std_logic;
signal \N__15493\ : std_logic;
signal \N__15490\ : std_logic;
signal \N__15487\ : std_logic;
signal \N__15484\ : std_logic;
signal \N__15483\ : std_logic;
signal \N__15482\ : std_logic;
signal \N__15481\ : std_logic;
signal \N__15480\ : std_logic;
signal \N__15477\ : std_logic;
signal \N__15476\ : std_logic;
signal \N__15475\ : std_logic;
signal \N__15474\ : std_logic;
signal \N__15473\ : std_logic;
signal \N__15472\ : std_logic;
signal \N__15467\ : std_logic;
signal \N__15462\ : std_logic;
signal \N__15459\ : std_logic;
signal \N__15456\ : std_logic;
signal \N__15451\ : std_logic;
signal \N__15446\ : std_logic;
signal \N__15443\ : std_logic;
signal \N__15440\ : std_logic;
signal \N__15435\ : std_logic;
signal \N__15434\ : std_logic;
signal \N__15429\ : std_logic;
signal \N__15424\ : std_logic;
signal \N__15421\ : std_logic;
signal \N__15418\ : std_logic;
signal \N__15409\ : std_logic;
signal \N__15406\ : std_logic;
signal \N__15403\ : std_logic;
signal \N__15400\ : std_logic;
signal \N__15397\ : std_logic;
signal \N__15394\ : std_logic;
signal \N__15391\ : std_logic;
signal \N__15388\ : std_logic;
signal \N__15385\ : std_logic;
signal \N__15384\ : std_logic;
signal \N__15381\ : std_logic;
signal \N__15378\ : std_logic;
signal \N__15377\ : std_logic;
signal \N__15374\ : std_logic;
signal \N__15371\ : std_logic;
signal \N__15368\ : std_logic;
signal \N__15363\ : std_logic;
signal \N__15358\ : std_logic;
signal \N__15357\ : std_logic;
signal \N__15352\ : std_logic;
signal \N__15349\ : std_logic;
signal \N__15346\ : std_logic;
signal \N__15343\ : std_logic;
signal \N__15340\ : std_logic;
signal \N__15337\ : std_logic;
signal \N__15336\ : std_logic;
signal \N__15333\ : std_logic;
signal \N__15330\ : std_logic;
signal \N__15327\ : std_logic;
signal \N__15324\ : std_logic;
signal \N__15321\ : std_logic;
signal \N__15320\ : std_logic;
signal \N__15317\ : std_logic;
signal \N__15314\ : std_logic;
signal \N__15311\ : std_logic;
signal \N__15304\ : std_logic;
signal \N__15301\ : std_logic;
signal \N__15298\ : std_logic;
signal \N__15297\ : std_logic;
signal \N__15294\ : std_logic;
signal \N__15291\ : std_logic;
signal \N__15286\ : std_logic;
signal \N__15283\ : std_logic;
signal \N__15280\ : std_logic;
signal \N__15279\ : std_logic;
signal \N__15276\ : std_logic;
signal \N__15273\ : std_logic;
signal \N__15268\ : std_logic;
signal \N__15265\ : std_logic;
signal \N__15262\ : std_logic;
signal \N__15259\ : std_logic;
signal \N__15256\ : std_logic;
signal \N__15253\ : std_logic;
signal \N__15250\ : std_logic;
signal \N__15247\ : std_logic;
signal \N__15244\ : std_logic;
signal \N__15241\ : std_logic;
signal \N__15238\ : std_logic;
signal \N__15235\ : std_logic;
signal \N__15232\ : std_logic;
signal \N__15229\ : std_logic;
signal \N__15226\ : std_logic;
signal \N__15223\ : std_logic;
signal \N__15220\ : std_logic;
signal \N__15217\ : std_logic;
signal \N__15214\ : std_logic;
signal \N__15211\ : std_logic;
signal \N__15208\ : std_logic;
signal \N__15205\ : std_logic;
signal \N__15202\ : std_logic;
signal \N__15199\ : std_logic;
signal \N__15196\ : std_logic;
signal \N__15193\ : std_logic;
signal \N__15192\ : std_logic;
signal \N__15189\ : std_logic;
signal \N__15186\ : std_logic;
signal \N__15181\ : std_logic;
signal \N__15178\ : std_logic;
signal \N__15175\ : std_logic;
signal \N__15172\ : std_logic;
signal \N__15169\ : std_logic;
signal \N__15166\ : std_logic;
signal \N__15163\ : std_logic;
signal \N__15160\ : std_logic;
signal \N__15157\ : std_logic;
signal \N__15154\ : std_logic;
signal \N__15151\ : std_logic;
signal \N__15148\ : std_logic;
signal \N__15145\ : std_logic;
signal \N__15142\ : std_logic;
signal \N__15139\ : std_logic;
signal \N__15136\ : std_logic;
signal \N__15133\ : std_logic;
signal \N__15130\ : std_logic;
signal \N__15127\ : std_logic;
signal \N__15126\ : std_logic;
signal \N__15121\ : std_logic;
signal \N__15118\ : std_logic;
signal \N__15117\ : std_logic;
signal \N__15112\ : std_logic;
signal \N__15111\ : std_logic;
signal \N__15110\ : std_logic;
signal \N__15109\ : std_logic;
signal \N__15108\ : std_logic;
signal \N__15107\ : std_logic;
signal \N__15104\ : std_logic;
signal \N__15099\ : std_logic;
signal \N__15096\ : std_logic;
signal \N__15091\ : std_logic;
signal \N__15088\ : std_logic;
signal \N__15081\ : std_logic;
signal \N__15076\ : std_logic;
signal \N__15073\ : std_logic;
signal \N__15072\ : std_logic;
signal \N__15067\ : std_logic;
signal \N__15064\ : std_logic;
signal \N__15061\ : std_logic;
signal \N__15060\ : std_logic;
signal \N__15059\ : std_logic;
signal \N__15056\ : std_logic;
signal \N__15055\ : std_logic;
signal \N__15050\ : std_logic;
signal \N__15047\ : std_logic;
signal \N__15044\ : std_logic;
signal \N__15041\ : std_logic;
signal \N__15040\ : std_logic;
signal \N__15039\ : std_logic;
signal \N__15038\ : std_logic;
signal \N__15035\ : std_logic;
signal \N__15032\ : std_logic;
signal \N__15029\ : std_logic;
signal \N__15022\ : std_logic;
signal \N__15013\ : std_logic;
signal \N__15010\ : std_logic;
signal \N__15007\ : std_logic;
signal \N__15004\ : std_logic;
signal \N__15001\ : std_logic;
signal \N__15000\ : std_logic;
signal \N__14995\ : std_logic;
signal \N__14992\ : std_logic;
signal \N__14989\ : std_logic;
signal \N__14986\ : std_logic;
signal \N__14983\ : std_logic;
signal \N__14980\ : std_logic;
signal \N__14977\ : std_logic;
signal \N__14974\ : std_logic;
signal \N__14971\ : std_logic;
signal \N__14968\ : std_logic;
signal \N__14965\ : std_logic;
signal \N__14962\ : std_logic;
signal \N__14959\ : std_logic;
signal \N__14956\ : std_logic;
signal \N__14953\ : std_logic;
signal \N__14950\ : std_logic;
signal \N__14947\ : std_logic;
signal \N__14944\ : std_logic;
signal \N__14941\ : std_logic;
signal \N__14938\ : std_logic;
signal \N__14935\ : std_logic;
signal \N__14932\ : std_logic;
signal \N__14929\ : std_logic;
signal \N__14926\ : std_logic;
signal \N__14923\ : std_logic;
signal \N__14920\ : std_logic;
signal \N__14919\ : std_logic;
signal \N__14918\ : std_logic;
signal \N__14917\ : std_logic;
signal \N__14910\ : std_logic;
signal \N__14909\ : std_logic;
signal \N__14908\ : std_logic;
signal \N__14907\ : std_logic;
signal \N__14906\ : std_logic;
signal \N__14903\ : std_logic;
signal \N__14900\ : std_logic;
signal \N__14899\ : std_logic;
signal \N__14898\ : std_logic;
signal \N__14891\ : std_logic;
signal \N__14888\ : std_logic;
signal \N__14885\ : std_logic;
signal \N__14882\ : std_logic;
signal \N__14877\ : std_logic;
signal \N__14874\ : std_logic;
signal \N__14863\ : std_logic;
signal \N__14860\ : std_logic;
signal \N__14857\ : std_logic;
signal \N__14854\ : std_logic;
signal \N__14851\ : std_logic;
signal \N__14848\ : std_logic;
signal \N__14845\ : std_logic;
signal \N__14842\ : std_logic;
signal \N__14841\ : std_logic;
signal \N__14840\ : std_logic;
signal \N__14839\ : std_logic;
signal \N__14838\ : std_logic;
signal \N__14837\ : std_logic;
signal \N__14836\ : std_logic;
signal \N__14835\ : std_logic;
signal \N__14826\ : std_logic;
signal \N__14817\ : std_logic;
signal \N__14812\ : std_logic;
signal \N__14811\ : std_logic;
signal \N__14810\ : std_logic;
signal \N__14809\ : std_logic;
signal \N__14808\ : std_logic;
signal \N__14805\ : std_logic;
signal \N__14804\ : std_logic;
signal \N__14803\ : std_logic;
signal \N__14800\ : std_logic;
signal \N__14797\ : std_logic;
signal \N__14796\ : std_logic;
signal \N__14795\ : std_logic;
signal \N__14786\ : std_logic;
signal \N__14777\ : std_logic;
signal \N__14774\ : std_logic;
signal \N__14767\ : std_logic;
signal \N__14766\ : std_logic;
signal \N__14765\ : std_logic;
signal \N__14764\ : std_logic;
signal \N__14763\ : std_logic;
signal \N__14762\ : std_logic;
signal \N__14761\ : std_logic;
signal \N__14758\ : std_logic;
signal \N__14755\ : std_logic;
signal \N__14754\ : std_logic;
signal \N__14751\ : std_logic;
signal \N__14742\ : std_logic;
signal \N__14733\ : std_logic;
signal \N__14728\ : std_logic;
signal \N__14727\ : std_logic;
signal \N__14724\ : std_logic;
signal \N__14721\ : std_logic;
signal \N__14720\ : std_logic;
signal \N__14719\ : std_logic;
signal \N__14718\ : std_logic;
signal \N__14717\ : std_logic;
signal \N__14716\ : std_logic;
signal \N__14715\ : std_logic;
signal \N__14706\ : std_logic;
signal \N__14697\ : std_logic;
signal \N__14692\ : std_logic;
signal \N__14689\ : std_logic;
signal \N__14686\ : std_logic;
signal \N__14683\ : std_logic;
signal \N__14680\ : std_logic;
signal \N__14677\ : std_logic;
signal \N__14674\ : std_logic;
signal \N__14671\ : std_logic;
signal \N__14668\ : std_logic;
signal \N__14665\ : std_logic;
signal \N__14662\ : std_logic;
signal \N__14659\ : std_logic;
signal \N__14656\ : std_logic;
signal \N__14653\ : std_logic;
signal \N__14650\ : std_logic;
signal \N__14647\ : std_logic;
signal \N__14644\ : std_logic;
signal \N__14641\ : std_logic;
signal \N__14640\ : std_logic;
signal \N__14635\ : std_logic;
signal \N__14632\ : std_logic;
signal \N__14629\ : std_logic;
signal \N__14626\ : std_logic;
signal \N__14623\ : std_logic;
signal \N__14620\ : std_logic;
signal \N__14617\ : std_logic;
signal \N__14614\ : std_logic;
signal \N__14611\ : std_logic;
signal \N__14608\ : std_logic;
signal \N__14605\ : std_logic;
signal \N__14602\ : std_logic;
signal \N__14599\ : std_logic;
signal \N__14596\ : std_logic;
signal \N__14593\ : std_logic;
signal \N__14590\ : std_logic;
signal \N__14589\ : std_logic;
signal \N__14586\ : std_logic;
signal \N__14585\ : std_logic;
signal \N__14578\ : std_logic;
signal \N__14575\ : std_logic;
signal \N__14572\ : std_logic;
signal \N__14569\ : std_logic;
signal \N__14566\ : std_logic;
signal \N__14563\ : std_logic;
signal \N__14560\ : std_logic;
signal \N__14557\ : std_logic;
signal \N__14554\ : std_logic;
signal \N__14551\ : std_logic;
signal \N__14548\ : std_logic;
signal \N__14545\ : std_logic;
signal \N__14542\ : std_logic;
signal \N__14539\ : std_logic;
signal \N__14536\ : std_logic;
signal \N__14533\ : std_logic;
signal \N__14530\ : std_logic;
signal \N__14527\ : std_logic;
signal \N__14524\ : std_logic;
signal \N__14521\ : std_logic;
signal \N__14518\ : std_logic;
signal \N__14515\ : std_logic;
signal \N__14512\ : std_logic;
signal \N__14509\ : std_logic;
signal \N__14508\ : std_logic;
signal \N__14505\ : std_logic;
signal \N__14502\ : std_logic;
signal \N__14501\ : std_logic;
signal \N__14500\ : std_logic;
signal \N__14497\ : std_logic;
signal \N__14494\ : std_logic;
signal \N__14491\ : std_logic;
signal \N__14488\ : std_logic;
signal \N__14483\ : std_logic;
signal \N__14480\ : std_logic;
signal \N__14477\ : std_logic;
signal \N__14474\ : std_logic;
signal \N__14467\ : std_logic;
signal \N__14464\ : std_logic;
signal \N__14461\ : std_logic;
signal \N__14458\ : std_logic;
signal \N__14455\ : std_logic;
signal \N__14452\ : std_logic;
signal \N__14449\ : std_logic;
signal \N__14446\ : std_logic;
signal \N__14443\ : std_logic;
signal \N__14440\ : std_logic;
signal \N__14437\ : std_logic;
signal \N__14434\ : std_logic;
signal \N__14431\ : std_logic;
signal \N__14428\ : std_logic;
signal \N__14427\ : std_logic;
signal \N__14424\ : std_logic;
signal \N__14421\ : std_logic;
signal \N__14416\ : std_logic;
signal \N__14415\ : std_logic;
signal \N__14414\ : std_logic;
signal \N__14413\ : std_logic;
signal \N__14410\ : std_logic;
signal \N__14407\ : std_logic;
signal \N__14402\ : std_logic;
signal \N__14395\ : std_logic;
signal \N__14392\ : std_logic;
signal \N__14389\ : std_logic;
signal \N__14386\ : std_logic;
signal \N__14383\ : std_logic;
signal \N__14380\ : std_logic;
signal \N__14379\ : std_logic;
signal \N__14376\ : std_logic;
signal \N__14375\ : std_logic;
signal \N__14372\ : std_logic;
signal \N__14367\ : std_logic;
signal \N__14362\ : std_logic;
signal \N__14361\ : std_logic;
signal \N__14358\ : std_logic;
signal \N__14353\ : std_logic;
signal \N__14350\ : std_logic;
signal \N__14347\ : std_logic;
signal \N__14344\ : std_logic;
signal \N__14341\ : std_logic;
signal \N__14338\ : std_logic;
signal \N__14335\ : std_logic;
signal \N__14332\ : std_logic;
signal \N__14329\ : std_logic;
signal \N__14328\ : std_logic;
signal \N__14323\ : std_logic;
signal \N__14320\ : std_logic;
signal \N__14317\ : std_logic;
signal \N__14314\ : std_logic;
signal \N__14313\ : std_logic;
signal \N__14308\ : std_logic;
signal \N__14305\ : std_logic;
signal \N__14304\ : std_logic;
signal \N__14299\ : std_logic;
signal \N__14296\ : std_logic;
signal \N__14293\ : std_logic;
signal \N__14292\ : std_logic;
signal \N__14289\ : std_logic;
signal \N__14286\ : std_logic;
signal \N__14283\ : std_logic;
signal \N__14278\ : std_logic;
signal \N__14275\ : std_logic;
signal \N__14272\ : std_logic;
signal \N__14269\ : std_logic;
signal \N__14268\ : std_logic;
signal \N__14265\ : std_logic;
signal \N__14262\ : std_logic;
signal \N__14259\ : std_logic;
signal \N__14256\ : std_logic;
signal \N__14253\ : std_logic;
signal \N__14250\ : std_logic;
signal \N__14247\ : std_logic;
signal \N__14242\ : std_logic;
signal \N__14239\ : std_logic;
signal \N__14236\ : std_logic;
signal \N__14233\ : std_logic;
signal \N__14230\ : std_logic;
signal \N__14227\ : std_logic;
signal \N__14224\ : std_logic;
signal \N__14223\ : std_logic;
signal \N__14222\ : std_logic;
signal \N__14219\ : std_logic;
signal \N__14214\ : std_logic;
signal \N__14209\ : std_logic;
signal \N__14206\ : std_logic;
signal \N__14205\ : std_logic;
signal \N__14202\ : std_logic;
signal \N__14199\ : std_logic;
signal \N__14194\ : std_logic;
signal \N__14191\ : std_logic;
signal \N__14188\ : std_logic;
signal \N__14185\ : std_logic;
signal \N__14182\ : std_logic;
signal \N__14179\ : std_logic;
signal \N__14176\ : std_logic;
signal \N__14175\ : std_logic;
signal \N__14172\ : std_logic;
signal \N__14169\ : std_logic;
signal \N__14164\ : std_logic;
signal \N__14161\ : std_logic;
signal \N__14160\ : std_logic;
signal \N__14157\ : std_logic;
signal \N__14156\ : std_logic;
signal \N__14153\ : std_logic;
signal \N__14150\ : std_logic;
signal \N__14147\ : std_logic;
signal \N__14140\ : std_logic;
signal \N__14137\ : std_logic;
signal \N__14134\ : std_logic;
signal \N__14131\ : std_logic;
signal \N__14128\ : std_logic;
signal \N__14125\ : std_logic;
signal \N__14122\ : std_logic;
signal \N__14119\ : std_logic;
signal \N__14116\ : std_logic;
signal \N__14113\ : std_logic;
signal \N__14110\ : std_logic;
signal \N__14107\ : std_logic;
signal \N__14104\ : std_logic;
signal \N__14101\ : std_logic;
signal \N__14098\ : std_logic;
signal \N__14097\ : std_logic;
signal \N__14096\ : std_logic;
signal \N__14095\ : std_logic;
signal \N__14092\ : std_logic;
signal \N__14089\ : std_logic;
signal \N__14088\ : std_logic;
signal \N__14087\ : std_logic;
signal \N__14084\ : std_logic;
signal \N__14083\ : std_logic;
signal \N__14080\ : std_logic;
signal \N__14077\ : std_logic;
signal \N__14064\ : std_logic;
signal \N__14059\ : std_logic;
signal \N__14056\ : std_logic;
signal \N__14053\ : std_logic;
signal \N__14050\ : std_logic;
signal \N__14047\ : std_logic;
signal \N__14044\ : std_logic;
signal \N__14041\ : std_logic;
signal \N__14038\ : std_logic;
signal \N__14035\ : std_logic;
signal \N__14034\ : std_logic;
signal \N__14033\ : std_logic;
signal \N__14026\ : std_logic;
signal \N__14025\ : std_logic;
signal \N__14022\ : std_logic;
signal \N__14019\ : std_logic;
signal \N__14016\ : std_logic;
signal \N__14011\ : std_logic;
signal \N__14008\ : std_logic;
signal \N__14007\ : std_logic;
signal \N__14004\ : std_logic;
signal \N__14001\ : std_logic;
signal \N__13998\ : std_logic;
signal \N__13995\ : std_logic;
signal \N__13992\ : std_logic;
signal \N__13987\ : std_logic;
signal \N__13984\ : std_logic;
signal \N__13981\ : std_logic;
signal \N__13978\ : std_logic;
signal \N__13975\ : std_logic;
signal \N__13974\ : std_logic;
signal \N__13971\ : std_logic;
signal \N__13968\ : std_logic;
signal \N__13965\ : std_logic;
signal \N__13962\ : std_logic;
signal \N__13957\ : std_logic;
signal \N__13954\ : std_logic;
signal \N__13951\ : std_logic;
signal \N__13948\ : std_logic;
signal \N__13945\ : std_logic;
signal \N__13942\ : std_logic;
signal \N__13939\ : std_logic;
signal \N__13938\ : std_logic;
signal \N__13935\ : std_logic;
signal \N__13932\ : std_logic;
signal \N__13929\ : std_logic;
signal \N__13926\ : std_logic;
signal \N__13921\ : std_logic;
signal \N__13920\ : std_logic;
signal \N__13917\ : std_logic;
signal \N__13914\ : std_logic;
signal \N__13909\ : std_logic;
signal \N__13906\ : std_logic;
signal \N__13903\ : std_logic;
signal \N__13900\ : std_logic;
signal \N__13897\ : std_logic;
signal \N__13896\ : std_logic;
signal \N__13893\ : std_logic;
signal \N__13890\ : std_logic;
signal \N__13887\ : std_logic;
signal \N__13884\ : std_logic;
signal \N__13881\ : std_logic;
signal \N__13878\ : std_logic;
signal \N__13873\ : std_logic;
signal \N__13870\ : std_logic;
signal \N__13867\ : std_logic;
signal \N__13864\ : std_logic;
signal \N__13863\ : std_logic;
signal \N__13862\ : std_logic;
signal \N__13859\ : std_logic;
signal \N__13854\ : std_logic;
signal \N__13851\ : std_logic;
signal \N__13848\ : std_logic;
signal \N__13845\ : std_logic;
signal \N__13842\ : std_logic;
signal \N__13837\ : std_logic;
signal \N__13834\ : std_logic;
signal \N__13831\ : std_logic;
signal \N__13830\ : std_logic;
signal \N__13829\ : std_logic;
signal \N__13824\ : std_logic;
signal \N__13821\ : std_logic;
signal \N__13818\ : std_logic;
signal \N__13815\ : std_logic;
signal \N__13812\ : std_logic;
signal \N__13809\ : std_logic;
signal \N__13804\ : std_logic;
signal \N__13801\ : std_logic;
signal \N__13798\ : std_logic;
signal \N__13795\ : std_logic;
signal \N__13792\ : std_logic;
signal \N__13789\ : std_logic;
signal \N__13786\ : std_logic;
signal \N__13783\ : std_logic;
signal \N__13780\ : std_logic;
signal \N__13777\ : std_logic;
signal \N__13774\ : std_logic;
signal \N__13771\ : std_logic;
signal \N__13768\ : std_logic;
signal \N__13765\ : std_logic;
signal \N__13762\ : std_logic;
signal \N__13759\ : std_logic;
signal \N__13756\ : std_logic;
signal \N__13753\ : std_logic;
signal \N__13750\ : std_logic;
signal \N__13747\ : std_logic;
signal \N__13744\ : std_logic;
signal \N__13741\ : std_logic;
signal \N__13738\ : std_logic;
signal \N__13735\ : std_logic;
signal \N__13732\ : std_logic;
signal \N__13729\ : std_logic;
signal \N__13726\ : std_logic;
signal \N__13725\ : std_logic;
signal \N__13722\ : std_logic;
signal \N__13719\ : std_logic;
signal \N__13714\ : std_logic;
signal \N__13711\ : std_logic;
signal \N__13708\ : std_logic;
signal \N__13705\ : std_logic;
signal \N__13702\ : std_logic;
signal \N__13699\ : std_logic;
signal \N__13696\ : std_logic;
signal \N__13693\ : std_logic;
signal \N__13692\ : std_logic;
signal \N__13689\ : std_logic;
signal \N__13688\ : std_logic;
signal \N__13685\ : std_logic;
signal \N__13684\ : std_logic;
signal \N__13681\ : std_logic;
signal \N__13674\ : std_logic;
signal \N__13669\ : std_logic;
signal \N__13666\ : std_logic;
signal \N__13663\ : std_logic;
signal \N__13662\ : std_logic;
signal \N__13659\ : std_logic;
signal \N__13656\ : std_logic;
signal \N__13655\ : std_logic;
signal \N__13654\ : std_logic;
signal \N__13651\ : std_logic;
signal \N__13648\ : std_logic;
signal \N__13643\ : std_logic;
signal \N__13636\ : std_logic;
signal \N__13633\ : std_logic;
signal \N__13630\ : std_logic;
signal \N__13627\ : std_logic;
signal \N__13626\ : std_logic;
signal \N__13625\ : std_logic;
signal \N__13624\ : std_logic;
signal \N__13623\ : std_logic;
signal \N__13620\ : std_logic;
signal \N__13615\ : std_logic;
signal \N__13610\ : std_logic;
signal \N__13603\ : std_logic;
signal \N__13600\ : std_logic;
signal \N__13597\ : std_logic;
signal \N__13594\ : std_logic;
signal \N__13593\ : std_logic;
signal \N__13590\ : std_logic;
signal \N__13589\ : std_logic;
signal \N__13586\ : std_logic;
signal \N__13585\ : std_logic;
signal \N__13584\ : std_logic;
signal \N__13583\ : std_logic;
signal \N__13580\ : std_logic;
signal \N__13573\ : std_logic;
signal \N__13568\ : std_logic;
signal \N__13561\ : std_logic;
signal \N__13558\ : std_logic;
signal \N__13557\ : std_logic;
signal \N__13556\ : std_logic;
signal \N__13553\ : std_logic;
signal \N__13550\ : std_logic;
signal \N__13547\ : std_logic;
signal \N__13544\ : std_logic;
signal \N__13539\ : std_logic;
signal \N__13534\ : std_logic;
signal \N__13531\ : std_logic;
signal \N__13528\ : std_logic;
signal \N__13525\ : std_logic;
signal \N__13522\ : std_logic;
signal \N__13519\ : std_logic;
signal \N__13516\ : std_logic;
signal \N__13513\ : std_logic;
signal \N__13510\ : std_logic;
signal \N__13507\ : std_logic;
signal \N__13504\ : std_logic;
signal \N__13501\ : std_logic;
signal \N__13498\ : std_logic;
signal \N__13495\ : std_logic;
signal \N__13492\ : std_logic;
signal \N__13489\ : std_logic;
signal \N__13486\ : std_logic;
signal \N__13483\ : std_logic;
signal \N__13480\ : std_logic;
signal \N__13477\ : std_logic;
signal \N__13474\ : std_logic;
signal \N__13471\ : std_logic;
signal \N__13468\ : std_logic;
signal \N__13467\ : std_logic;
signal \N__13466\ : std_logic;
signal \N__13463\ : std_logic;
signal \N__13460\ : std_logic;
signal \N__13457\ : std_logic;
signal \N__13454\ : std_logic;
signal \N__13451\ : std_logic;
signal \N__13450\ : std_logic;
signal \N__13447\ : std_logic;
signal \N__13444\ : std_logic;
signal \N__13441\ : std_logic;
signal \N__13438\ : std_logic;
signal \N__13435\ : std_logic;
signal \N__13426\ : std_logic;
signal \N__13425\ : std_logic;
signal \N__13422\ : std_logic;
signal \N__13419\ : std_logic;
signal \N__13416\ : std_logic;
signal \N__13411\ : std_logic;
signal \N__13408\ : std_logic;
signal \N__13407\ : std_logic;
signal \N__13402\ : std_logic;
signal \N__13399\ : std_logic;
signal \N__13396\ : std_logic;
signal \N__13393\ : std_logic;
signal \N__13390\ : std_logic;
signal \N__13387\ : std_logic;
signal \N__13384\ : std_logic;
signal \N__13383\ : std_logic;
signal \N__13380\ : std_logic;
signal \N__13377\ : std_logic;
signal \N__13372\ : std_logic;
signal \N__13369\ : std_logic;
signal \N__13366\ : std_logic;
signal \N__13363\ : std_logic;
signal \N__13360\ : std_logic;
signal \N__13357\ : std_logic;
signal \N__13356\ : std_logic;
signal \N__13355\ : std_logic;
signal \N__13352\ : std_logic;
signal \N__13349\ : std_logic;
signal \N__13346\ : std_logic;
signal \N__13339\ : std_logic;
signal \N__13336\ : std_logic;
signal \N__13333\ : std_logic;
signal \N__13330\ : std_logic;
signal \N__13329\ : std_logic;
signal \N__13326\ : std_logic;
signal \N__13321\ : std_logic;
signal \N__13318\ : std_logic;
signal \N__13315\ : std_logic;
signal \N__13312\ : std_logic;
signal \N__13309\ : std_logic;
signal \N__13308\ : std_logic;
signal \N__13307\ : std_logic;
signal \N__13300\ : std_logic;
signal \N__13297\ : std_logic;
signal \N__13296\ : std_logic;
signal \N__13293\ : std_logic;
signal \N__13292\ : std_logic;
signal \N__13285\ : std_logic;
signal \N__13282\ : std_logic;
signal \N__13279\ : std_logic;
signal \N__13276\ : std_logic;
signal \N__13273\ : std_logic;
signal \N__13270\ : std_logic;
signal \N__13267\ : std_logic;
signal \N__13264\ : std_logic;
signal \N__13261\ : std_logic;
signal \N__13258\ : std_logic;
signal \N__13255\ : std_logic;
signal \N__13252\ : std_logic;
signal \N__13249\ : std_logic;
signal \N__13246\ : std_logic;
signal \N__13243\ : std_logic;
signal \N__13240\ : std_logic;
signal \N__13237\ : std_logic;
signal \N__13234\ : std_logic;
signal \N__13233\ : std_logic;
signal \N__13230\ : std_logic;
signal \N__13227\ : std_logic;
signal \N__13224\ : std_logic;
signal \N__13223\ : std_logic;
signal \N__13220\ : std_logic;
signal \N__13217\ : std_logic;
signal \N__13216\ : std_logic;
signal \N__13213\ : std_logic;
signal \N__13210\ : std_logic;
signal \N__13207\ : std_logic;
signal \N__13204\ : std_logic;
signal \N__13195\ : std_logic;
signal \N__13192\ : std_logic;
signal \N__13191\ : std_logic;
signal \N__13186\ : std_logic;
signal \N__13183\ : std_logic;
signal \N__13182\ : std_logic;
signal \N__13177\ : std_logic;
signal \N__13174\ : std_logic;
signal \N__13171\ : std_logic;
signal \N__13168\ : std_logic;
signal \N__13167\ : std_logic;
signal \N__13162\ : std_logic;
signal \N__13159\ : std_logic;
signal \N__13156\ : std_logic;
signal \N__13153\ : std_logic;
signal \N__13150\ : std_logic;
signal \N__13147\ : std_logic;
signal \N__13144\ : std_logic;
signal \N__13141\ : std_logic;
signal \N__13138\ : std_logic;
signal \N__13135\ : std_logic;
signal \N__13132\ : std_logic;
signal \N__13129\ : std_logic;
signal \N__13126\ : std_logic;
signal \N__13123\ : std_logic;
signal \N__13120\ : std_logic;
signal \N__13117\ : std_logic;
signal \N__13116\ : std_logic;
signal \N__13115\ : std_logic;
signal \N__13114\ : std_logic;
signal \N__13113\ : std_logic;
signal \N__13106\ : std_logic;
signal \N__13103\ : std_logic;
signal \N__13100\ : std_logic;
signal \N__13097\ : std_logic;
signal \N__13090\ : std_logic;
signal \N__13089\ : std_logic;
signal \N__13088\ : std_logic;
signal \N__13085\ : std_logic;
signal \N__13080\ : std_logic;
signal \N__13079\ : std_logic;
signal \N__13078\ : std_logic;
signal \N__13077\ : std_logic;
signal \N__13074\ : std_logic;
signal \N__13071\ : std_logic;
signal \N__13066\ : std_logic;
signal \N__13063\ : std_logic;
signal \N__13060\ : std_logic;
signal \N__13057\ : std_logic;
signal \N__13048\ : std_logic;
signal \N__13045\ : std_logic;
signal \N__13044\ : std_logic;
signal \N__13039\ : std_logic;
signal \N__13036\ : std_logic;
signal \N__13033\ : std_logic;
signal \N__13030\ : std_logic;
signal \N__13027\ : std_logic;
signal \N__13024\ : std_logic;
signal \N__13023\ : std_logic;
signal \N__13018\ : std_logic;
signal \N__13015\ : std_logic;
signal \N__13012\ : std_logic;
signal \N__13011\ : std_logic;
signal \N__13008\ : std_logic;
signal \N__13007\ : std_logic;
signal \N__13004\ : std_logic;
signal \N__13001\ : std_logic;
signal \N__12998\ : std_logic;
signal \N__12995\ : std_logic;
signal \N__12990\ : std_logic;
signal \N__12989\ : std_logic;
signal \N__12988\ : std_logic;
signal \N__12987\ : std_logic;
signal \N__12986\ : std_logic;
signal \N__12985\ : std_logic;
signal \N__12984\ : std_logic;
signal \N__12983\ : std_logic;
signal \N__12982\ : std_logic;
signal \N__12981\ : std_logic;
signal \N__12978\ : std_logic;
signal \N__12975\ : std_logic;
signal \N__12968\ : std_logic;
signal \N__12963\ : std_logic;
signal \N__12954\ : std_logic;
signal \N__12951\ : std_logic;
signal \N__12940\ : std_logic;
signal \N__12939\ : std_logic;
signal \N__12938\ : std_logic;
signal \N__12935\ : std_logic;
signal \N__12932\ : std_logic;
signal \N__12929\ : std_logic;
signal \N__12926\ : std_logic;
signal \N__12919\ : std_logic;
signal \N__12916\ : std_logic;
signal \N__12915\ : std_logic;
signal \N__12912\ : std_logic;
signal \N__12909\ : std_logic;
signal \N__12906\ : std_logic;
signal \N__12903\ : std_logic;
signal \N__12900\ : std_logic;
signal \N__12897\ : std_logic;
signal \N__12892\ : std_logic;
signal \N__12889\ : std_logic;
signal \N__12886\ : std_logic;
signal \N__12883\ : std_logic;
signal \N__12880\ : std_logic;
signal \N__12877\ : std_logic;
signal \N__12874\ : std_logic;
signal \N__12871\ : std_logic;
signal \N__12870\ : std_logic;
signal \N__12865\ : std_logic;
signal \N__12862\ : std_logic;
signal \N__12859\ : std_logic;
signal \N__12856\ : std_logic;
signal \N__12853\ : std_logic;
signal \N__12850\ : std_logic;
signal \N__12847\ : std_logic;
signal \N__12844\ : std_logic;
signal \N__12841\ : std_logic;
signal \N__12838\ : std_logic;
signal \N__12835\ : std_logic;
signal \N__12832\ : std_logic;
signal \N__12831\ : std_logic;
signal \N__12830\ : std_logic;
signal \N__12827\ : std_logic;
signal \N__12826\ : std_logic;
signal \N__12825\ : std_logic;
signal \N__12820\ : std_logic;
signal \N__12819\ : std_logic;
signal \N__12818\ : std_logic;
signal \N__12817\ : std_logic;
signal \N__12816\ : std_logic;
signal \N__12815\ : std_logic;
signal \N__12814\ : std_logic;
signal \N__12813\ : std_logic;
signal \N__12812\ : std_logic;
signal \N__12811\ : std_logic;
signal \N__12808\ : std_logic;
signal \N__12803\ : std_logic;
signal \N__12800\ : std_logic;
signal \N__12799\ : std_logic;
signal \N__12798\ : std_logic;
signal \N__12781\ : std_logic;
signal \N__12778\ : std_logic;
signal \N__12771\ : std_logic;
signal \N__12766\ : std_logic;
signal \N__12757\ : std_logic;
signal \N__12754\ : std_logic;
signal \N__12751\ : std_logic;
signal \N__12748\ : std_logic;
signal \N__12745\ : std_logic;
signal \N__12742\ : std_logic;
signal \N__12739\ : std_logic;
signal \N__12736\ : std_logic;
signal \N__12733\ : std_logic;
signal \N__12730\ : std_logic;
signal \N__12729\ : std_logic;
signal \N__12726\ : std_logic;
signal \N__12723\ : std_logic;
signal \N__12720\ : std_logic;
signal \N__12717\ : std_logic;
signal \N__12712\ : std_logic;
signal \N__12709\ : std_logic;
signal \N__12706\ : std_logic;
signal \N__12703\ : std_logic;
signal \N__12700\ : std_logic;
signal \N__12697\ : std_logic;
signal \N__12694\ : std_logic;
signal \N__12691\ : std_logic;
signal \N__12688\ : std_logic;
signal \N__12685\ : std_logic;
signal \N__12682\ : std_logic;
signal \N__12679\ : std_logic;
signal \N__12676\ : std_logic;
signal \N__12673\ : std_logic;
signal \N__12670\ : std_logic;
signal \N__12667\ : std_logic;
signal \N__12666\ : std_logic;
signal \N__12661\ : std_logic;
signal \N__12658\ : std_logic;
signal \N__12655\ : std_logic;
signal \N__12652\ : std_logic;
signal \N__12649\ : std_logic;
signal \N__12646\ : std_logic;
signal \N__12643\ : std_logic;
signal \N__12640\ : std_logic;
signal \N__12637\ : std_logic;
signal \N__12634\ : std_logic;
signal \N__12631\ : std_logic;
signal \N__12628\ : std_logic;
signal \N__12625\ : std_logic;
signal \N__12622\ : std_logic;
signal \N__12619\ : std_logic;
signal \N__12616\ : std_logic;
signal \N__12613\ : std_logic;
signal \N__12610\ : std_logic;
signal \N__12609\ : std_logic;
signal \N__12606\ : std_logic;
signal \N__12603\ : std_logic;
signal \N__12600\ : std_logic;
signal \N__12595\ : std_logic;
signal \N__12592\ : std_logic;
signal \N__12589\ : std_logic;
signal \N__12586\ : std_logic;
signal \N__12583\ : std_logic;
signal \N__12580\ : std_logic;
signal \N__12577\ : std_logic;
signal \N__12574\ : std_logic;
signal \N__12571\ : std_logic;
signal \N__12568\ : std_logic;
signal \N__12565\ : std_logic;
signal \N__12562\ : std_logic;
signal \N__12559\ : std_logic;
signal \N__12556\ : std_logic;
signal \N__12553\ : std_logic;
signal \N__12550\ : std_logic;
signal \N__12547\ : std_logic;
signal \N__12544\ : std_logic;
signal \N__12541\ : std_logic;
signal \N__12538\ : std_logic;
signal \N__12535\ : std_logic;
signal \N__12532\ : std_logic;
signal \N__12529\ : std_logic;
signal \N__12526\ : std_logic;
signal \N__12525\ : std_logic;
signal \N__12524\ : std_logic;
signal \N__12523\ : std_logic;
signal \N__12514\ : std_logic;
signal \N__12513\ : std_logic;
signal \N__12512\ : std_logic;
signal \N__12509\ : std_logic;
signal \N__12506\ : std_logic;
signal \N__12503\ : std_logic;
signal \N__12498\ : std_logic;
signal \N__12493\ : std_logic;
signal \N__12490\ : std_logic;
signal \N__12487\ : std_logic;
signal \N__12484\ : std_logic;
signal \N__12481\ : std_logic;
signal \N__12480\ : std_logic;
signal \N__12475\ : std_logic;
signal \N__12474\ : std_logic;
signal \N__12473\ : std_logic;
signal \N__12470\ : std_logic;
signal \N__12467\ : std_logic;
signal \N__12464\ : std_logic;
signal \N__12461\ : std_logic;
signal \N__12458\ : std_logic;
signal \N__12451\ : std_logic;
signal \N__12450\ : std_logic;
signal \N__12449\ : std_logic;
signal \N__12446\ : std_logic;
signal \N__12441\ : std_logic;
signal \N__12438\ : std_logic;
signal \N__12433\ : std_logic;
signal \N__12430\ : std_logic;
signal \N__12427\ : std_logic;
signal \N__12426\ : std_logic;
signal \N__12423\ : std_logic;
signal \N__12420\ : std_logic;
signal \N__12417\ : std_logic;
signal \N__12412\ : std_logic;
signal \N__12411\ : std_logic;
signal \N__12406\ : std_logic;
signal \N__12403\ : std_logic;
signal \N__12402\ : std_logic;
signal \N__12401\ : std_logic;
signal \N__12400\ : std_logic;
signal \N__12397\ : std_logic;
signal \N__12394\ : std_logic;
signal \N__12389\ : std_logic;
signal \N__12382\ : std_logic;
signal \N__12379\ : std_logic;
signal \N__12376\ : std_logic;
signal \N__12375\ : std_logic;
signal \N__12374\ : std_logic;
signal \N__12373\ : std_logic;
signal \N__12370\ : std_logic;
signal \N__12367\ : std_logic;
signal \N__12364\ : std_logic;
signal \N__12361\ : std_logic;
signal \N__12358\ : std_logic;
signal \N__12355\ : std_logic;
signal \N__12346\ : std_logic;
signal \N__12345\ : std_logic;
signal \N__12344\ : std_logic;
signal \N__12343\ : std_logic;
signal \N__12342\ : std_logic;
signal \N__12331\ : std_logic;
signal \N__12328\ : std_logic;
signal \N__12325\ : std_logic;
signal \N__12322\ : std_logic;
signal \N__12319\ : std_logic;
signal \N__12316\ : std_logic;
signal \N__12313\ : std_logic;
signal \N__12310\ : std_logic;
signal \N__12307\ : std_logic;
signal \N__12304\ : std_logic;
signal \N__12301\ : std_logic;
signal \N__12298\ : std_logic;
signal \N__12295\ : std_logic;
signal \N__12292\ : std_logic;
signal \N__12289\ : std_logic;
signal \N__12286\ : std_logic;
signal \N__12283\ : std_logic;
signal \N__12280\ : std_logic;
signal \N__12277\ : std_logic;
signal \N__12274\ : std_logic;
signal \N__12271\ : std_logic;
signal \N__12268\ : std_logic;
signal \N__12265\ : std_logic;
signal \N__12262\ : std_logic;
signal \N__12259\ : std_logic;
signal \N__12256\ : std_logic;
signal \N__12253\ : std_logic;
signal \N__12250\ : std_logic;
signal \N__12247\ : std_logic;
signal \N__12244\ : std_logic;
signal \N__12241\ : std_logic;
signal \N__12238\ : std_logic;
signal \N__12235\ : std_logic;
signal \N__12232\ : std_logic;
signal \N__12229\ : std_logic;
signal \N__12226\ : std_logic;
signal \N__12223\ : std_logic;
signal \N__12220\ : std_logic;
signal \N__12217\ : std_logic;
signal \N__12214\ : std_logic;
signal \N__12211\ : std_logic;
signal \N__12208\ : std_logic;
signal \N__12205\ : std_logic;
signal \N__12202\ : std_logic;
signal \N__12201\ : std_logic;
signal \N__12200\ : std_logic;
signal \N__12199\ : std_logic;
signal \N__12198\ : std_logic;
signal \N__12187\ : std_logic;
signal \N__12184\ : std_logic;
signal \N__12183\ : std_logic;
signal \N__12182\ : std_logic;
signal \N__12181\ : std_logic;
signal \N__12178\ : std_logic;
signal \N__12177\ : std_logic;
signal \N__12172\ : std_logic;
signal \N__12165\ : std_logic;
signal \N__12160\ : std_logic;
signal \N__12159\ : std_logic;
signal \N__12158\ : std_logic;
signal \N__12155\ : std_logic;
signal \N__12148\ : std_logic;
signal \N__12145\ : std_logic;
signal \N__12142\ : std_logic;
signal \N__12139\ : std_logic;
signal \N__12136\ : std_logic;
signal \N__12133\ : std_logic;
signal \N__12130\ : std_logic;
signal \N__12127\ : std_logic;
signal \N__12126\ : std_logic;
signal \N__12125\ : std_logic;
signal \N__12124\ : std_logic;
signal \N__12123\ : std_logic;
signal \N__12112\ : std_logic;
signal \N__12109\ : std_logic;
signal \N__12108\ : std_logic;
signal \N__12107\ : std_logic;
signal \N__12100\ : std_logic;
signal \N__12097\ : std_logic;
signal \N__12094\ : std_logic;
signal \N__12091\ : std_logic;
signal \N__12088\ : std_logic;
signal \N__12085\ : std_logic;
signal \N__12082\ : std_logic;
signal \N__12079\ : std_logic;
signal \N__12078\ : std_logic;
signal \N__12077\ : std_logic;
signal \N__12074\ : std_logic;
signal \N__12071\ : std_logic;
signal \N__12068\ : std_logic;
signal \N__12065\ : std_logic;
signal \N__12058\ : std_logic;
signal \N__12057\ : std_logic;
signal \N__12056\ : std_logic;
signal \N__12053\ : std_logic;
signal \N__12048\ : std_logic;
signal \N__12043\ : std_logic;
signal \N__12042\ : std_logic;
signal \N__12039\ : std_logic;
signal \N__12036\ : std_logic;
signal \N__12031\ : std_logic;
signal \N__12028\ : std_logic;
signal \N__12025\ : std_logic;
signal \N__12024\ : std_logic;
signal \N__12023\ : std_logic;
signal \N__12022\ : std_logic;
signal \N__12019\ : std_logic;
signal \N__12012\ : std_logic;
signal \N__12007\ : std_logic;
signal \N__12006\ : std_logic;
signal \N__12005\ : std_logic;
signal \N__12000\ : std_logic;
signal \N__11997\ : std_logic;
signal \N__11992\ : std_logic;
signal \N__11989\ : std_logic;
signal \N__11986\ : std_logic;
signal \N__11983\ : std_logic;
signal \N__11980\ : std_logic;
signal \N__11977\ : std_logic;
signal \N__11974\ : std_logic;
signal \N__11971\ : std_logic;
signal \N__11968\ : std_logic;
signal \N__11965\ : std_logic;
signal \N__11962\ : std_logic;
signal \N__11959\ : std_logic;
signal \N__11956\ : std_logic;
signal \N__11953\ : std_logic;
signal \N__11950\ : std_logic;
signal \N__11947\ : std_logic;
signal \N__11944\ : std_logic;
signal \N__11941\ : std_logic;
signal \N__11938\ : std_logic;
signal \N__11935\ : std_logic;
signal \N__11932\ : std_logic;
signal \N__11929\ : std_logic;
signal \N__11926\ : std_logic;
signal \N__11923\ : std_logic;
signal \N__11920\ : std_logic;
signal \N__11917\ : std_logic;
signal \N__11914\ : std_logic;
signal \N__11911\ : std_logic;
signal \N__11908\ : std_logic;
signal \N__11905\ : std_logic;
signal \N__11902\ : std_logic;
signal \N__11899\ : std_logic;
signal \N__11896\ : std_logic;
signal \N__11893\ : std_logic;
signal \N__11890\ : std_logic;
signal \N__11887\ : std_logic;
signal \N__11884\ : std_logic;
signal \N__11881\ : std_logic;
signal \N__11878\ : std_logic;
signal \N__11875\ : std_logic;
signal \N__11872\ : std_logic;
signal \N__11871\ : std_logic;
signal \N__11870\ : std_logic;
signal \N__11869\ : std_logic;
signal \N__11868\ : std_logic;
signal \N__11857\ : std_logic;
signal \N__11854\ : std_logic;
signal \N__11853\ : std_logic;
signal \N__11852\ : std_logic;
signal \N__11849\ : std_logic;
signal \N__11846\ : std_logic;
signal \N__11839\ : std_logic;
signal \N__11836\ : std_logic;
signal \N__11835\ : std_logic;
signal \N__11834\ : std_logic;
signal \N__11831\ : std_logic;
signal \N__11830\ : std_logic;
signal \N__11823\ : std_logic;
signal \N__11820\ : std_logic;
signal \N__11815\ : std_logic;
signal \N__11814\ : std_logic;
signal \N__11811\ : std_logic;
signal \N__11808\ : std_logic;
signal \N__11803\ : std_logic;
signal \N__11802\ : std_logic;
signal \N__11801\ : std_logic;
signal \N__11798\ : std_logic;
signal \N__11793\ : std_logic;
signal \N__11790\ : std_logic;
signal \N__11785\ : std_logic;
signal \N__11782\ : std_logic;
signal \N__11779\ : std_logic;
signal \N__11776\ : std_logic;
signal \N__11773\ : std_logic;
signal \N__11770\ : std_logic;
signal \N__11767\ : std_logic;
signal \N__11764\ : std_logic;
signal \N__11761\ : std_logic;
signal \N__11758\ : std_logic;
signal \N__11755\ : std_logic;
signal \N__11752\ : std_logic;
signal \N__11749\ : std_logic;
signal \N__11746\ : std_logic;
signal \N__11743\ : std_logic;
signal \N__11740\ : std_logic;
signal \N__11737\ : std_logic;
signal \N__11736\ : std_logic;
signal \N__11735\ : std_logic;
signal \N__11734\ : std_logic;
signal \N__11733\ : std_logic;
signal \N__11732\ : std_logic;
signal \N__11729\ : std_logic;
signal \N__11726\ : std_logic;
signal \N__11725\ : std_logic;
signal \N__11724\ : std_logic;
signal \N__11723\ : std_logic;
signal \N__11720\ : std_logic;
signal \N__11717\ : std_logic;
signal \N__11716\ : std_logic;
signal \N__11709\ : std_logic;
signal \N__11706\ : std_logic;
signal \N__11699\ : std_logic;
signal \N__11692\ : std_logic;
signal \N__11683\ : std_logic;
signal \N__11682\ : std_logic;
signal \N__11681\ : std_logic;
signal \N__11676\ : std_logic;
signal \N__11673\ : std_logic;
signal \N__11670\ : std_logic;
signal \N__11665\ : std_logic;
signal \N__11662\ : std_logic;
signal \N__11661\ : std_logic;
signal \N__11660\ : std_logic;
signal \N__11659\ : std_logic;
signal \N__11654\ : std_logic;
signal \N__11649\ : std_logic;
signal \N__11644\ : std_logic;
signal \N__11641\ : std_logic;
signal \N__11640\ : std_logic;
signal \N__11639\ : std_logic;
signal \N__11638\ : std_logic;
signal \N__11637\ : std_logic;
signal \N__11630\ : std_logic;
signal \N__11625\ : std_logic;
signal \N__11620\ : std_logic;
signal \N__11617\ : std_logic;
signal \N__11616\ : std_logic;
signal \N__11615\ : std_logic;
signal \N__11608\ : std_logic;
signal \N__11605\ : std_logic;
signal \N__11604\ : std_logic;
signal \N__11603\ : std_logic;
signal \N__11600\ : std_logic;
signal \N__11593\ : std_logic;
signal \N__11590\ : std_logic;
signal \N__11589\ : std_logic;
signal \N__11588\ : std_logic;
signal \N__11583\ : std_logic;
signal \N__11580\ : std_logic;
signal \N__11575\ : std_logic;
signal \N__11572\ : std_logic;
signal \N__11569\ : std_logic;
signal \N__11566\ : std_logic;
signal \N__11565\ : std_logic;
signal \N__11564\ : std_logic;
signal \N__11563\ : std_logic;
signal \N__11560\ : std_logic;
signal \N__11557\ : std_logic;
signal \N__11554\ : std_logic;
signal \N__11551\ : std_logic;
signal \N__11550\ : std_logic;
signal \N__11547\ : std_logic;
signal \N__11544\ : std_logic;
signal \N__11537\ : std_logic;
signal \N__11530\ : std_logic;
signal \N__11527\ : std_logic;
signal \N__11526\ : std_logic;
signal \N__11525\ : std_logic;
signal \N__11524\ : std_logic;
signal \N__11523\ : std_logic;
signal \N__11520\ : std_logic;
signal \N__11519\ : std_logic;
signal \N__11518\ : std_logic;
signal \N__11517\ : std_logic;
signal \N__11516\ : std_logic;
signal \N__11513\ : std_logic;
signal \N__11506\ : std_logic;
signal \N__11503\ : std_logic;
signal \N__11494\ : std_logic;
signal \N__11491\ : std_logic;
signal \N__11482\ : std_logic;
signal \N__11481\ : std_logic;
signal \N__11480\ : std_logic;
signal \N__11477\ : std_logic;
signal \N__11474\ : std_logic;
signal \N__11471\ : std_logic;
signal \N__11468\ : std_logic;
signal \N__11465\ : std_logic;
signal \N__11458\ : std_logic;
signal \N__11457\ : std_logic;
signal \N__11456\ : std_logic;
signal \N__11455\ : std_logic;
signal \N__11452\ : std_logic;
signal \N__11445\ : std_logic;
signal \N__11442\ : std_logic;
signal \N__11437\ : std_logic;
signal \N__11434\ : std_logic;
signal \N__11431\ : std_logic;
signal \N__11428\ : std_logic;
signal \N__11425\ : std_logic;
signal \N__11422\ : std_logic;
signal \N__11419\ : std_logic;
signal \N__11418\ : std_logic;
signal \N__11415\ : std_logic;
signal \N__11414\ : std_logic;
signal \N__11409\ : std_logic;
signal \N__11406\ : std_logic;
signal \N__11401\ : std_logic;
signal \N__11398\ : std_logic;
signal \N__11397\ : std_logic;
signal \N__11396\ : std_logic;
signal \N__11395\ : std_logic;
signal \N__11386\ : std_logic;
signal \N__11383\ : std_logic;
signal \N__11382\ : std_logic;
signal \N__11381\ : std_logic;
signal \N__11380\ : std_logic;
signal \N__11375\ : std_logic;
signal \N__11370\ : std_logic;
signal \N__11365\ : std_logic;
signal \N__11362\ : std_logic;
signal \N__11361\ : std_logic;
signal \N__11360\ : std_logic;
signal \N__11357\ : std_logic;
signal \N__11352\ : std_logic;
signal \N__11347\ : std_logic;
signal \N__11346\ : std_logic;
signal \N__11345\ : std_logic;
signal \N__11344\ : std_logic;
signal \N__11341\ : std_logic;
signal \N__11336\ : std_logic;
signal \N__11331\ : std_logic;
signal \N__11326\ : std_logic;
signal \N__11325\ : std_logic;
signal \N__11324\ : std_logic;
signal \N__11323\ : std_logic;
signal \N__11322\ : std_logic;
signal \N__11321\ : std_logic;
signal \N__11318\ : std_logic;
signal \N__11313\ : std_logic;
signal \N__11306\ : std_logic;
signal \N__11299\ : std_logic;
signal \N__11296\ : std_logic;
signal \N__11293\ : std_logic;
signal \N__11290\ : std_logic;
signal \N__11287\ : std_logic;
signal \N__11284\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11278\ : std_logic;
signal \N__11275\ : std_logic;
signal \N__11272\ : std_logic;
signal \N__11269\ : std_logic;
signal \N__11268\ : std_logic;
signal \N__11267\ : std_logic;
signal \N__11266\ : std_logic;
signal \N__11259\ : std_logic;
signal \N__11256\ : std_logic;
signal \N__11251\ : std_logic;
signal \N__11248\ : std_logic;
signal \N__11245\ : std_logic;
signal \N__11242\ : std_logic;
signal \N__11239\ : std_logic;
signal \N__11236\ : std_logic;
signal \N__11233\ : std_logic;
signal \N__11230\ : std_logic;
signal \N__11227\ : std_logic;
signal \N__11224\ : std_logic;
signal \N__11221\ : std_logic;
signal \N__11218\ : std_logic;
signal \N__11215\ : std_logic;
signal \N__11212\ : std_logic;
signal \N__11209\ : std_logic;
signal \N__11206\ : std_logic;
signal \N__11203\ : std_logic;
signal \N__11200\ : std_logic;
signal \N__11197\ : std_logic;
signal \N__11196\ : std_logic;
signal \N__11191\ : std_logic;
signal \N__11188\ : std_logic;
signal \N__11185\ : std_logic;
signal \N__11184\ : std_logic;
signal \N__11179\ : std_logic;
signal \N__11176\ : std_logic;
signal \N__11175\ : std_logic;
signal \N__11172\ : std_logic;
signal \N__11169\ : std_logic;
signal \N__11166\ : std_logic;
signal \N__11161\ : std_logic;
signal \N__11160\ : std_logic;
signal \N__11155\ : std_logic;
signal \N__11152\ : std_logic;
signal \N__11151\ : std_logic;
signal \N__11146\ : std_logic;
signal \N__11143\ : std_logic;
signal \N__11140\ : std_logic;
signal \N__11139\ : std_logic;
signal \N__11136\ : std_logic;
signal \N__11135\ : std_logic;
signal \N__11132\ : std_logic;
signal \N__11127\ : std_logic;
signal \N__11122\ : std_logic;
signal \N__11121\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11119\ : std_logic;
signal \N__11114\ : std_logic;
signal \N__11109\ : std_logic;
signal \N__11104\ : std_logic;
signal \N__11101\ : std_logic;
signal \N__11098\ : std_logic;
signal \N__11095\ : std_logic;
signal \N__11092\ : std_logic;
signal \N__11089\ : std_logic;
signal \N__11086\ : std_logic;
signal \N__11083\ : std_logic;
signal \N__11080\ : std_logic;
signal \N__11077\ : std_logic;
signal \N__11076\ : std_logic;
signal \N__11073\ : std_logic;
signal \N__11070\ : std_logic;
signal \N__11065\ : std_logic;
signal \N__11064\ : std_logic;
signal \N__11061\ : std_logic;
signal \N__11058\ : std_logic;
signal \N__11055\ : std_logic;
signal \N__11050\ : std_logic;
signal \N__11047\ : std_logic;
signal \N__11046\ : std_logic;
signal \N__11043\ : std_logic;
signal \N__11040\ : std_logic;
signal \N__11035\ : std_logic;
signal \N__11032\ : std_logic;
signal \N__11029\ : std_logic;
signal \N__11028\ : std_logic;
signal \N__11027\ : std_logic;
signal \N__11024\ : std_logic;
signal \N__11023\ : std_logic;
signal \N__11022\ : std_logic;
signal \N__11011\ : std_logic;
signal \N__11008\ : std_logic;
signal \N__11005\ : std_logic;
signal \N__11002\ : std_logic;
signal \N__10999\ : std_logic;
signal \N__10996\ : std_logic;
signal \N__10993\ : std_logic;
signal \N__10990\ : std_logic;
signal \N__10987\ : std_logic;
signal \N__10984\ : std_logic;
signal \N__10981\ : std_logic;
signal \N__10978\ : std_logic;
signal \N__10975\ : std_logic;
signal \N__10974\ : std_logic;
signal \N__10969\ : std_logic;
signal \N__10966\ : std_logic;
signal \N__10965\ : std_logic;
signal \N__10964\ : std_logic;
signal \N__10957\ : std_logic;
signal \N__10954\ : std_logic;
signal \N__10951\ : std_logic;
signal \N__10948\ : std_logic;
signal \N__10945\ : std_logic;
signal \N__10942\ : std_logic;
signal \N__10939\ : std_logic;
signal \N__10936\ : std_logic;
signal \N__10933\ : std_logic;
signal \N__10930\ : std_logic;
signal \latticehx1k_pll_inst.clk\ : std_logic;
signal clk_in_c : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \uu0.un187_ci_1_cascade_\ : std_logic;
signal \uu0.un165_ci_0\ : std_logic;
signal \uu0.l_countZ0Z_13\ : std_logic;
signal \uu0.l_countZ0Z_12\ : std_logic;
signal \uu0.un4_l_count_0_8_cascade_\ : std_logic;
signal \uu0.l_countZ0Z_0\ : std_logic;
signal \uu0.un44_ci\ : std_logic;
signal \uu0.un44_ci_cascade_\ : std_logic;
signal \bfn_1_4_0_\ : std_logic;
signal \buart.Z_tx.un1_bitcount_cry_0\ : std_logic;
signal \buart.Z_tx.bitcount_RNIVE1P1_0Z0Z_3\ : std_logic;
signal \buart.Z_tx.un1_bitcount_cry_1\ : std_logic;
signal \buart.Z_tx.un1_bitcount_cry_2\ : std_logic;
signal \buart.Z_tx.bitcount_RNIVE1P1Z0Z_3\ : std_logic;
signal \buart.Z_tx.un1_bitcount_axb_3\ : std_logic;
signal \buart.Z_tx.un1_bitcount_cry_0_0_c_RNOZ0\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_1\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_3\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_2\ : std_logic;
signal \buart.Z_tx.uart_busy_0_i_cascade_\ : std_logic;
signal \bfn_1_6_0_\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_1\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_2\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_3\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_4\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_5\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_5\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_4\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_6\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_3\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_2\ : std_logic;
signal \buart.Z_tx.Z_baudgen.ser_clk_4_cascade_\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_1\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_0\ : std_logic;
signal \Lab_UT.dictrl.N_17_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g0_i_4_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_19\ : std_logic;
signal \Lab_UT.dictrl.N_8_2\ : std_logic;
signal \Lab_UT.dictrl.N_8_2_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g0_i_a8_0_1\ : std_logic;
signal \Lab_UT.dictrl.N_1605_1\ : std_logic;
signal \Lab_UT.dictrl.currState_0_ret_28_RNOZ0Z_4_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_1605_0\ : std_logic;
signal \Lab_UT.dictrl.N_5_0\ : std_logic;
signal \Lab_UT.dictrl.g1_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g0_i_o4_4_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g0_i_o4_4_cascade_\ : std_logic;
signal \uart_RXD\ : std_logic;
signal \uu0.l_countZ0Z_2\ : std_logic;
signal \uu0.un4_l_count_14_cascade_\ : std_logic;
signal \uu0.un4_l_count_13\ : std_logic;
signal \uu0.un4_l_count_18_cascade_\ : std_logic;
signal \uu0.un4_l_count_0_cascade_\ : std_logic;
signal \uu0.un143_ci_0\ : std_logic;
signal \uu0.l_countZ0Z_11\ : std_logic;
signal \uu0.l_countZ0Z_10\ : std_logic;
signal \uu0.un154_ci_9\ : std_logic;
signal \uu0.un154_ci_9_cascade_\ : std_logic;
signal \uu0.un4_l_count_0_8\ : std_logic;
signal \uu0.l_countZ0Z_14\ : std_logic;
signal \uu0.l_countZ0Z_8\ : std_logic;
signal \uu0.un110_ci\ : std_logic;
signal \uu0.un198_ci_2\ : std_logic;
signal \uu0.un110_ci_cascade_\ : std_logic;
signal \uu0.l_countZ0Z_16\ : std_logic;
signal \uu0.un220_ci_cascade_\ : std_logic;
signal \uu0.l_countZ0Z_9\ : std_logic;
signal \uu0.l_countZ0Z_7\ : std_logic;
signal \uu0.l_countZ0Z_17\ : std_logic;
signal \uu0.l_countZ0Z_3\ : std_logic;
signal \uu0.un4_l_count_12\ : std_logic;
signal \buart.Z_tx.uart_busy_0_i\ : std_logic;
signal \buart.Z_tx.ser_clk\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_0\ : std_logic;
signal \uu0.l_precountZ0Z_2\ : std_logic;
signal \uu0.l_precountZ0Z_1\ : std_logic;
signal \uu0.l_precountZ0Z_3\ : std_logic;
signal \uu0.l_countZ0Z_1\ : std_logic;
signal \uu0.l_countZ0Z_18\ : std_logic;
signal \uu0.l_countZ0Z_15\ : std_logic;
signal \uu0.un4_l_count_11_cascade_\ : std_logic;
signal \uu0.un4_l_count_16\ : std_logic;
signal \uu2.r_data_wire_0\ : std_logic;
signal \uu2.r_data_wire_1\ : std_logic;
signal \uu2.r_data_wire_2\ : std_logic;
signal \uu2.r_data_wire_3\ : std_logic;
signal \uu2.r_data_wire_4\ : std_logic;
signal \uu2.r_data_wire_5\ : std_logic;
signal \uu2.r_data_wire_6\ : std_logic;
signal \uu2.r_data_wire_7\ : std_logic;
signal \INVuu2.r_data_reg_0C_net\ : std_logic;
signal vbuf_tx_data_0 : std_logic;
signal \buart.Z_tx.shifterZ0Z_1\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_0\ : std_logic;
signal o_serial_data_c : std_logic;
signal vbuf_tx_data_1 : std_logic;
signal \buart.Z_tx.shifterZ0Z_2\ : std_logic;
signal vbuf_tx_data_2 : std_logic;
signal \buart.Z_tx.shifterZ0Z_3\ : std_logic;
signal vbuf_tx_data_3 : std_logic;
signal \buart.Z_tx.shifterZ0Z_4\ : std_logic;
signal vbuf_tx_data_4 : std_logic;
signal \buart.Z_tx.shifterZ0Z_5\ : std_logic;
signal vbuf_tx_data_5 : std_logic;
signal \buart.Z_tx.shifterZ0Z_6\ : std_logic;
signal \INVuu2.vram_rd_clk_det_0C_net\ : std_logic;
signal \uu2.un1_l_count_1_3_cascade_\ : std_logic;
signal \uu2.un1_l_count_1_3\ : std_logic;
signal \uu2.un1_l_count_2_0_cascade_\ : std_logic;
signal \uu2.l_countZ0Z_2\ : std_logic;
signal \uu2.l_countZ0Z_3\ : std_logic;
signal \uu2.un306_ci_cascade_\ : std_logic;
signal \uu2.un350_ci_cascade_\ : std_logic;
signal \uu2.un1_l_count_1_2_0\ : std_logic;
signal \uu2.un350_ci\ : std_logic;
signal \uu2.l_countZ0Z_8\ : std_logic;
signal \uu2.l_countZ0Z_5\ : std_logic;
signal \uu2.vbuf_count.un328_ci_3\ : std_logic;
signal \uu2.vbuf_count.un328_ci_3_cascade_\ : std_logic;
signal \uu2.un306_ci\ : std_logic;
signal \uu2.l_countZ0Z_7\ : std_logic;
signal \uu2.l_countZ0Z_6\ : std_logic;
signal \uu2.l_countZ0Z_4\ : std_logic;
signal \uu2.l_countZ0Z_9\ : std_logic;
signal \uu2.un1_l_count_2_2\ : std_logic;
signal \Lab_UT.dictrl.N_8_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_20_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_9_1\ : std_logic;
signal \Lab_UT.dictrl.G_30_0_a7_4_1\ : std_logic;
signal \Lab_UT.dictrl.G_30_0_a7_1_2\ : std_logic;
signal \Lab_UT.dictrl.N_31_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_23_1\ : std_logic;
signal \Lab_UT.dictrl.G_30_0_2_cascade_\ : std_logic;
signal \Lab_UT.dictrl.nextStateZ0Z_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.G_30_0_a7_2_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.G_30_0_0\ : std_logic;
signal \Lab_UT.dictrl.G_30_0_a7_0_0\ : std_logic;
signal \Lab_UT.dictrl.N_30_0\ : std_logic;
signal \Lab_UT.dictrl.i8_mux_0_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.i7_mux_0\ : std_logic;
signal \Lab_UT.dictrl.N_12\ : std_logic;
signal \Lab_UT.dictrl.G_30_0_a7_2\ : std_logic;
signal \Lab_UT.dictrl.N_11_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_5_0_0\ : std_logic;
signal \Lab_UT.dictrl.g0_4_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_8_0_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_4\ : std_logic;
signal \Lab_UT.dictrl.currState_i_5_2\ : std_logic;
signal \Lab_UT.dictrl.G_19_0_a7_4_10_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_21_cascade_\ : std_logic;
signal \Lab_UT.dictrl.G_19_0_a7_2_0\ : std_logic;
signal \Lab_UT.dictrl.G_19_0_0\ : std_logic;
signal \Lab_UT.dictrl.G_19_0_a7_3_2\ : std_logic;
signal \G_19_0_a7_4_8\ : std_logic;
signal \G_19_0_a7_4_1\ : std_logic;
signal \uu0.l_precountZ0Z_0\ : std_logic;
signal \uu0.un99_ci_0\ : std_logic;
signal \uu0.l_countZ0Z_4\ : std_logic;
signal \uu0.l_countZ0Z_5\ : std_logic;
signal \uu0.un88_ci_3\ : std_logic;
signal \uu0.un66_ci\ : std_logic;
signal \uu0.un88_ci_3_cascade_\ : std_logic;
signal \uu0.l_countZ0Z_6\ : std_logic;
signal \uu0.un11_l_count_i_g\ : std_logic;
signal \uu2.mem0.w_addr_8\ : std_logic;
signal \uu2.vram_rd_clk_detZ0Z_1\ : std_logic;
signal \uu2.vram_rd_clk_detZ0Z_0\ : std_logic;
signal \uu2.vram_rd_clk_det_RNI95711Z0Z_1\ : std_logic;
signal \uu2.mem0.w_data_4\ : std_logic;
signal \uu2.mem0.w_data_5\ : std_logic;
signal \uu2.N_37\ : std_logic;
signal \uu2.N_37_cascade_\ : std_logic;
signal \uu2.mem0.w_data_3\ : std_logic;
signal \uu2.mem0.w_data_1\ : std_logic;
signal \uu2.N_51_cascade_\ : std_logic;
signal \uu2.N_34\ : std_logic;
signal \uu2.N_34_cascade_\ : std_logic;
signal \uu2.mem0.w_data_0\ : std_logic;
signal \uu2.bitmap_pmux_sn_m15_0_ns_1_cascade_\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_65\ : std_logic;
signal \uu2.bitmap_pmux_sn_m24_0_ns_1_cascade_\ : std_logic;
signal \uu2.bitmap_pmux_sn_i5_mux_cascade_\ : std_logic;
signal \uu2.bitmap_pmux_sn_i7_mux_0\ : std_logic;
signal \uu2.bitmap_pmux_29_0_cascade_\ : std_logic;
signal \uu2.bitmap_pmux\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_36\ : std_logic;
signal vbuf_tx_data_6 : std_logic;
signal \buart.Z_tx.shifterZ0Z_7\ : std_logic;
signal vbuf_tx_data_rdy : std_logic;
signal vbuf_tx_data_7 : std_logic;
signal \buart.Z_tx.shifterZ0Z_8\ : std_logic;
signal \buart.Z_tx.un1_uart_wr_i_0_i\ : std_logic;
signal \uu0.un11_l_count_i\ : std_logic;
signal \uu2.mem0.w_addr_7\ : std_logic;
signal \uu2.mem0.w_addr_1\ : std_logic;
signal \uu2.w_data_displaying_2_i_a2_i_a3_1_0\ : std_logic;
signal \uu0.un4_l_count_0\ : std_logic;
signal \uu2.un1_l_count_2_0\ : std_logic;
signal \uu0.delay_lineZ0Z_0\ : std_logic;
signal \uu0.delay_lineZ0Z_1\ : std_logic;
signal \uu2.l_countZ0Z_1\ : std_logic;
signal \uu2.l_countZ0Z_0\ : std_logic;
signal \uu2.un284_ci\ : std_logic;
signal \Lab_UT.dictrl.N_9_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_21_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g0_0_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_1611_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_23_0\ : std_logic;
signal \Lab_UT.dictrl.N_8_3\ : std_logic;
signal \Lab_UT.dictrl.G_28_0_a5_1\ : std_logic;
signal \Lab_UT.dictrl.N_19_0\ : std_logic;
signal \Lab_UT.dictrl.N_8_3_cascade_\ : std_logic;
signal \Lab_UT.dictrl.currState_2_0_rep2_RNIBGCIZ0Z9_cascade_\ : std_logic;
signal \Lab_UT.dictrl.G_28_0_0\ : std_logic;
signal \Lab_UT.dictrl.currState_2_0_rep2_RNIKH8PZ0Z2\ : std_logic;
signal \shifter_RNIS6CF1_5\ : std_logic;
signal \Lab_UT.dictrl.m21_rn_1_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.m21_rn_0\ : std_logic;
signal \Lab_UT.dictrl.g1_0_1\ : std_logic;
signal \Lab_UT.dictrl.N_7_1\ : std_logic;
signal \Lab_UT.dictrl.nextState_0_1\ : std_logic;
signal \Lab_UT.dictrl.N_20_cascade_\ : std_logic;
signal \Lab_UT.dictrl.decoder.g0Z0Z_5_cascade_\ : std_logic;
signal \Lab_UT.dictrl.decoder.g0Z0Z_1\ : std_logic;
signal \Lab_UT.dictrl.N_36_1_cascade_\ : std_logic;
signal \G_28_0_a5_0_4_cascade_\ : std_logic;
signal \shifter_RNI1D8L1_4\ : std_logic;
signal \bfn_4_16_0_\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_1\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_2\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_3\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_4\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_5\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_2\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_1\ : std_logic;
signal \uu2.trig_rd_is_det_cascade_\ : std_logic;
signal \uu2.trig_rd_detZ0Z_1\ : std_logic;
signal \uu2.vram_rd_clkZ0\ : std_logic;
signal \uu2.un1_l_count_1_0\ : std_logic;
signal \uu2.trig_rd_detZ0Z_0\ : std_logic;
signal \uu2.vbuf_raddr.un448_ci_0\ : std_logic;
signal \uu2.vbuf_raddr.un426_ci_3_cascade_\ : std_logic;
signal \uu2.r_addrZ0Z_8\ : std_logic;
signal \uu2.vbuf_raddr.un426_ci_3\ : std_logic;
signal \uu2.r_addrZ0Z_7\ : std_logic;
signal \uu2.un404_ci_0_cascade_\ : std_logic;
signal \uu2.r_addrZ0Z_6\ : std_logic;
signal \uu2.r_addrZ0Z_2\ : std_logic;
signal \uu2.r_addrZ0Z_1\ : std_logic;
signal \uu2.r_addrZ0Z_0\ : std_logic;
signal \uu2.r_addrZ0Z_3\ : std_logic;
signal \uu2.trig_rd_is_det_0\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_42\ : std_logic;
signal \uu2.bitmap_pmux_26_bm_1_cascade_\ : std_logic;
signal \uu2.N_161\ : std_logic;
signal \uu2.N_400_cascade_\ : std_logic;
signal \uu2.N_409\ : std_logic;
signal \uu2.bitmap_RNI1PH82Z0Z_34\ : std_logic;
signal \uu2.N_404\ : std_logic;
signal \uu2.bitmapZ0Z_290\ : std_logic;
signal \uu2.bitmapZ0Z_40\ : std_logic;
signal \uu2.bitmapZ0Z_296\ : std_logic;
signal \INVuu2.bitmap_290C_net\ : std_logic;
signal \uu2.bitmap_pmux_25_am_1_cascade_\ : std_logic;
signal \uu2.bitmapZ0Z_197\ : std_logic;
signal \uu2.bitmapZ0Z_66\ : std_logic;
signal \INVuu2.bitmap_197C_net\ : std_logic;
signal \uu2.bitmap_RNI2JA82Z0Z_212_cascade_\ : std_logic;
signal \uu2.N_31_i\ : std_logic;
signal \uu2.bitmap_RNIM7D32Z0Z_69\ : std_logic;
signal \uu2.bitmap_pmux_27_ns_1_cascade_\ : std_logic;
signal \uu2.N_407\ : std_logic;
signal \Lab_UT.segmentUQ_0_0_cascade_\ : std_logic;
signal \Lab_UT.N_65_0_cascade_\ : std_logic;
signal \Lab_UT.segment_1_0_6\ : std_logic;
signal \Lab_UT.N_76_0_cascade_\ : std_logic;
signal \INVuu2.bitmap_72C_net\ : std_logic;
signal \uu2.bitmapZ0Z_72\ : std_logic;
signal \uu2.bitmapZ0Z_200\ : std_logic;
signal \uu2.bitmap_RNIOS152Z0Z_72\ : std_logic;
signal \Lab_UT.dictrl.currState_ret_RNI7FNUZ0\ : std_logic;
signal \Lab_UT.Mone_at_0_cascade_\ : std_logic;
signal \Lab_UT.N_77_0\ : std_logic;
signal \Lab_UT.dictrl.N_23\ : std_logic;
signal \Lab_UT.dictrl.N_23_cascade_\ : std_logic;
signal \Lab_UT.dictrl.nextState_RNIA8EV3Z0Z_1\ : std_logic;
signal \Lab_UT.dictrl.N_10\ : std_logic;
signal \Lab_UT.dictrl.N_12_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.G_28_0_a5_2_1\ : std_logic;
signal \Lab_UT.dictrl.dicLdAMtensZ0\ : std_logic;
signal \Lab_UT.dictrl.dicLdAMtens_rst\ : std_logic;
signal \Lab_UT.dictrl.r_dicLdMtens16_1\ : std_logic;
signal \Lab_UT.dictrl.g0_10_0_N_4L6_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.r_dicLdMtens17_1\ : std_logic;
signal \Lab_UT.dictrl.r_dicLdMtens22_2\ : std_logic;
signal \Lab_UT.dictrl.N_34_cascade_\ : std_logic;
signal \Lab_UT.dictrl.currState_2_RNI0P25DZ0Z_1\ : std_logic;
signal \Lab_UT.dictrl.m15_bm_cascade_\ : std_logic;
signal \Lab_UT.dictrl.nextState_0_0\ : std_logic;
signal \Lab_UT.dictrl.N_7_0\ : std_logic;
signal \Lab_UT.dictrl.N_1609_1\ : std_logic;
signal \Lab_UT.dictrl.N_38\ : std_logic;
signal \Lab_UT.dictrl.currState_ret_5_RNOZ0Z_0\ : std_logic;
signal \Lab_UT.dictrl.N_23_0_0\ : std_logic;
signal \Lab_UT.dictrl.N_13_0_0\ : std_logic;
signal \Lab_UT.dictrl.N_14_0_0_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_1609_0_0\ : std_logic;
signal \Lab_UT.dictrl.N_8\ : std_logic;
signal \Lab_UT.dictrl.N_7\ : std_logic;
signal \Lab_UT.dictrl.N_9_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g0_6\ : std_logic;
signal \Lab_UT.dictrl.N_6_0\ : std_logic;
signal \Lab_UT.dictrl.N_9\ : std_logic;
signal \Lab_UT.dictrl.m15_am\ : std_logic;
signal \Lab_UT.dictrl.N_20_1\ : std_logic;
signal \Lab_UT.dictrl.currState_0_rep1\ : std_logic;
signal \buart.Z_rx.bitcount_fast_es_RNIAJ1GZ0Z_3_cascade_\ : std_logic;
signal \bu_rx_data_rdy_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_5_0_1\ : std_logic;
signal \Lab_UT.dictrl.g0_3_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g0_1_0_0\ : std_logic;
signal bu_rx_data_fast_0 : std_logic;
signal \Lab_UT.dictrl.de_num_1_2\ : std_logic;
signal bu_rx_data_fast_7 : std_logic;
signal \Lab_UT.dictrl.decoder.g0_5_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.de_cr_0_0\ : std_logic;
signal \Lab_UT.dictrl.decoder.g0_6_0\ : std_logic;
signal bu_rx_data_fast_6 : std_logic;
signal \Lab_UT.dictrl.decoder.g0Z0Z_4\ : std_logic;
signal bu_rx_data_fast_4 : std_logic;
signal bu_rx_data_fast_5 : std_logic;
signal \buart.Z_rx.hhZ0Z_0\ : std_logic;
signal \Lab_UT.dictrl.decoder.g0Z0Z_7_cascade_\ : std_logic;
signal \Lab_UT.dictrl.currState_fast_0\ : std_logic;
signal \Lab_UT.dictrl.g1_4_1_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.de_littleA_0\ : std_logic;
signal \Lab_UT.dictrl.g1_4_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_17_0_0\ : std_logic;
signal \Lab_UT.dictrl.decoder.g0_5_1\ : std_logic;
signal \Lab_UT.dictrl.m7_sx\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_3\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_0\ : std_logic;
signal \buart.Z_rx.Z_baudgen.ser_clk_3\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO\ : std_logic;
signal \buart.Z_rx.ser_clk_cascade_\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_4\ : std_logic;
signal \resetGen.reset_count_2_0_4_cascade_\ : std_logic;
signal \uu2.mem0.w_addr_2\ : std_logic;
signal \uu2.mem0.w_addr_4\ : std_logic;
signal \uu2.mem0.w_addr_5\ : std_logic;
signal \uu2.mem0.w_addr_6\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_20\ : std_logic;
signal \uu2.bitmapZ0Z_168\ : std_logic;
signal \uu2.N_17_cascade_\ : std_logic;
signal \uu2.bitmap_RNIELSJ2Z0Z_111\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_54_mux\ : std_logic;
signal \uu2.bitmapZ0Z_111\ : std_logic;
signal \INVuu2.bitmap_111C_net\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_33\ : std_logic;
signal \uu2.N_39_cascade_\ : std_logic;
signal \uu2.N_48\ : std_logic;
signal \INVuu2.w_addr_displaying_nesr_3C_net\ : std_logic;
signal \uu2.bitmap_pmux_24_am_1\ : std_logic;
signal \uu2.bitmapZ0Z_87\ : std_logic;
signal \uu2.N_386_cascade_\ : std_logic;
signal \uu2.w_addr_displaying_nesr_RNI1JET2Z0Z_7_cascade_\ : std_logic;
signal \uu2.bitmapZ0Z_314\ : std_logic;
signal \uu2.bitmap_pmux_23_ns_1\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_15\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_2\ : std_logic;
signal \INVuu2.bitmap_87C_net\ : std_logic;
signal \Lab_UT.L3_segment3_0_i_1_0\ : std_logic;
signal \Lab_UT.L3_segment3_0_i_1_3\ : std_logic;
signal \Lab_UT.L3_segment3_1_2_cascade_\ : std_logic;
signal \Lab_UT.Mone_at_0\ : std_logic;
signal \Lab_UT.Mone_at_3\ : std_logic;
signal \Lab_UT.Mone_at_2\ : std_logic;
signal \Lab_UT.Mone_at_1\ : std_logic;
signal \Lab_UT.L3_segment3_1_1_cascade_\ : std_logic;
signal \uu2.bitmapZ0Z_203\ : std_logic;
signal \uu2.bitmapZ0Z_75\ : std_logic;
signal \uu2.bitmap_pmux_24_bm_1\ : std_logic;
signal \INVuu2.bitmap_203C_net\ : std_logic;
signal \Lab_UT.N_76_cascade_\ : std_logic;
signal \uu2.bitmapZ0Z_194\ : std_logic;
signal \Lab_UT.L3_segment4_1_1_cascade_\ : std_logic;
signal \uu2.bitmapZ0Z_69\ : std_logic;
signal \Lab_UT.L3_segment4_1_0\ : std_logic;
signal \uu2.bitmapZ0Z_34\ : std_logic;
signal \Lab_UT.segment_1_6_cascade_\ : std_logic;
signal \uu2.bitmapZ0Z_162\ : std_logic;
signal \INVuu2.bitmap_194C_net\ : std_logic;
signal \Lab_UT.dictrl.N_1614_0\ : std_logic;
signal \Lab_UT.dictrl.N_26\ : std_logic;
signal \Lab_UT.dictrl.un1_currState_6\ : std_logic;
signal \Lab_UT.dictrl.r_enableZ0Z1\ : std_logic;
signal \Lab_UT.dictrl.enableSeg3\ : std_logic;
signal \Lab_UT.dictrl.r_enableZ0Z3\ : std_logic;
signal \Lab_UT.dictrl.enableSeg4\ : std_logic;
signal \Lab_UT.dictrl.un1_currState_7\ : std_logic;
signal \Lab_UT.dictrl.r_enableZ0Z4\ : std_logic;
signal \Lab_UT.dictrl.N_1605_1_0\ : std_logic;
signal \Lab_UT.dictrl.N_36_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.nextStateZ0Z_3_cascade_\ : std_logic;
signal \Lab_UT.dictrl.r_dicLdMtens21_1\ : std_logic;
signal \Lab_UT.dictrl.N_18\ : std_logic;
signal \Lab_UT.dictrl.N_33\ : std_logic;
signal \Lab_UT.dictrl.N_1607_0_0\ : std_logic;
signal \Lab_UT.dictrl.N_10_0_0\ : std_logic;
signal \Lab_UT.dictrl.g1\ : std_logic;
signal \Lab_UT.dictrl.g2_cascade_\ : std_logic;
signal \Lab_UT.dictrl.nextState_RNO_9Z0Z_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g0_i_a4_1\ : std_logic;
signal \Lab_UT.dictrl.nextState_RNO_4Z0Z_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.nextState_RNO_3Z0Z_1\ : std_logic;
signal \Lab_UT.dictrl.g0_i_o4_5\ : std_logic;
signal \Lab_UT.dictrl.N_11\ : std_logic;
signal \Lab_UT.dictrl.N_18_0\ : std_logic;
signal \Lab_UT.dictrl.g1_3_0\ : std_logic;
signal \Lab_UT.dictrl.N_13_0\ : std_logic;
signal \Lab_UT.dictrl.g1_4_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_14\ : std_logic;
signal \Lab_UT.dictrl.r_dicLdMtens20_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_6ctr\ : std_logic;
signal \Lab_UT.dictrl.r_dicLdMtens22_2_reti\ : std_logic;
signal \Lab_UT.dictrl.N_7_1_0\ : std_logic;
signal \Lab_UT.dictrl.r_dicLdMtens22_2_reti_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g0_0_3\ : std_logic;
signal \Lab_UT.dictrl.N_10ctr\ : std_logic;
signal \Lab_UT.dictrl.r_dicLdMtens22_4_0\ : std_logic;
signal \N_7\ : std_logic;
signal \Lab_UT.dictrl.N_20\ : std_logic;
signal \Lab_UT.dictrl.de_littleA\ : std_logic;
signal \Lab_UT_dictrl_decoder_de_cr_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_30\ : std_logic;
signal \Lab_UT.dictrl.N_41_mux\ : std_logic;
signal \Lab_UT.dictrl.N_34\ : std_logic;
signal \Lab_UT.dictrl.N_31_cascade_\ : std_logic;
signal \Lab_UT.dictrl.nextState_0_2\ : std_logic;
signal \Lab_UT.dictrl.currState_0_ret_29_RNIDFRSEEZ0\ : std_logic;
signal \buart__rx_bitcount_fast_2\ : std_logic;
signal \buart__rx_bitcount_fast_4\ : std_logic;
signal \buart__rx_bitcount_fast_3\ : std_logic;
signal \Lab_UT.dictrl.decoder.g0_6_1\ : std_logic;
signal \buart.Z_rx.un1_sample_0_cascade_\ : std_logic;
signal \buart.Z_rx.sample\ : std_logic;
signal \buart.Z_rx.idle_0_cascade_\ : std_logic;
signal \buart.Z_rx.idle\ : std_logic;
signal \buart.Z_rx.ser_clk\ : std_logic;
signal \buart.Z_rx.idle_cascade_\ : std_logic;
signal \buart.Z_rx.N_27_0_i\ : std_logic;
signal \buart.Z_rx.startbit\ : std_logic;
signal \buart.Z_rx.bitcounte_0_0\ : std_logic;
signal \buart__rx_bitcount_0\ : std_logic;
signal \bfn_6_16_0_\ : std_logic;
signal \buart__rx_bitcount_1\ : std_logic;
signal \buart.Z_rx.bitcount_cry_0_THRU_CO\ : std_logic;
signal \buart.Z_rx.bitcount_cry_0\ : std_logic;
signal \buart.Z_rx.bitcount_cry_1_THRU_CO\ : std_logic;
signal \buart.Z_rx.bitcount_cry_1\ : std_logic;
signal \buart.Z_rx.bitcount_cry_2_THRU_CO\ : std_logic;
signal \buart.Z_rx.bitcount_cry_2\ : std_logic;
signal \buart.Z_rx.bitcount_cry_3\ : std_logic;
signal \buart.Z_rx.bitcount_cry_3_THRU_CO\ : std_logic;
signal \Lab_UT.uu0.l_countZ0Z_13\ : std_logic;
signal \Lab_UT.uu0.un143_ci_0_cascade_\ : std_logic;
signal \Lab_UT.uu0.un154_ci_9_cascade_\ : std_logic;
signal \Lab_UT.uu0.l_countZ0Z_12\ : std_logic;
signal \Lab_UT.uu0.un165_ci_0\ : std_logic;
signal \uu2.un3_w_addr_user_4_cascade_\ : std_logic;
signal \uu2.un3_w_addr_user_5\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_3\ : std_logic;
signal \uu2.mem0.w_addr_3\ : std_logic;
signal \uu2.vbuf_w_addr_user.un448_ci_0_cascade_\ : std_logic;
signal \uu2.w_addr_userZ0Z_8\ : std_logic;
signal \uu2.w_addr_userZ0Z_7\ : std_logic;
signal \INVuu2.w_addr_user_nesr_3C_net\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_1\ : std_logic;
signal \uu2.N_39\ : std_logic;
signal \INVuu2.w_addr_displaying_8C_net\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_5\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_4\ : std_logic;
signal \uu2.N_41\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_6\ : std_logic;
signal \uu2.N_41_cascade_\ : std_logic;
signal \uu2.N_43\ : std_logic;
signal \uu2.N_40\ : std_logic;
signal \uu2.N_43_cascade_\ : std_logic;
signal \uu2.w_addr_displaying_RNIFCPV4Z0Z_8\ : std_logic;
signal \uu2.w_addr_displaying_RNIFCPV4Z0Z_8_cascade_\ : std_logic;
signal \uu2.N_36_0\ : std_logic;
signal \Lab_UT.L3_segment2_1_1\ : std_logic;
signal \Lab_UT.L3_segment2_0_i_1_3_cascade_\ : std_logic;
signal \Lab_UT.L3_segment2_1_2_cascade_\ : std_logic;
signal \uu2.bitmapZ0Z_215\ : std_logic;
signal \Lab_UT.L3_segment2_0_i_1_0_cascade_\ : std_logic;
signal \INVuu2.bitmap_308C_net\ : std_logic;
signal \uu2.bitmapZ0Z_52\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_8\ : std_logic;
signal \uu2.bitmapZ0Z_308\ : std_logic;
signal \uu2.N_158\ : std_logic;
signal \Lab_UT.segmentUQ_0_0_1_cascade_\ : std_logic;
signal \Lab_UT.N_65_2_cascade_\ : std_logic;
signal \Lab_UT.segment_1_2_6\ : std_logic;
signal \uu2.bitmapZ0Z_186\ : std_logic;
signal \Lab_UT.N_76_2_cascade_\ : std_logic;
signal \INVuu2.bitmap_90C_net\ : std_logic;
signal \uu2.bitmapZ0Z_90\ : std_logic;
signal \uu2.bitmapZ0Z_218\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_7\ : std_logic;
signal \Lab_UT.N_76_1_cascade_\ : std_logic;
signal \uu2.bitmapZ0Z_212\ : std_logic;
signal \Lab_UT.N_65_1_cascade_\ : std_logic;
signal \Lab_UT.segment_1_1_6\ : std_logic;
signal \uu2.bitmapZ0Z_180\ : std_logic;
signal \Lab_UT.N_77_1\ : std_logic;
signal \uu2.bitmapZ0Z_84\ : std_logic;
signal \INVuu2.bitmap_212C_net\ : std_logic;
signal \Lab_UT.L3_segment4_0_i_1_5\ : std_logic;
signal \Lab_UT.N_65\ : std_logic;
signal \Lab_UT.Mten_at_3_cascade_\ : std_logic;
signal \Lab_UT.segment_1_3\ : std_logic;
signal \Lab_UT.N_69_0\ : std_logic;
signal \Lab_UT.N_69_0_cascade_\ : std_logic;
signal \Lab_UT.N_92\ : std_logic;
signal \Lab_UT.N_67_0\ : std_logic;
signal \Lab_UT.N_91\ : std_logic;
signal \Lab_UT.N_83\ : std_logic;
signal \Lab_UT.Mten_at_0\ : std_logic;
signal \Lab_UT.Mten_at_3\ : std_logic;
signal \Lab_UT.Mten_at_0_cascade_\ : std_logic;
signal \Lab_UT.N_77\ : std_logic;
signal \Lab_UT.Mten_at_1\ : std_logic;
signal \Lab_UT.dictrl.g0_13_1\ : std_logic;
signal \Lab_UT.dictrl.g0_1\ : std_logic;
signal \Lab_UT.dictrl.g0_i_o4_0_0\ : std_logic;
signal \Lab_UT.dictrl.currState_0_ret_20and_1_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.de_cr\ : std_logic;
signal \Lab_UT.dictrl.N_13\ : std_logic;
signal \Lab_UT.dictrl.N_17_0\ : std_logic;
signal \Lab_UT.dictrl.N_13_cascade_\ : std_logic;
signal \Lab_UT.dictrl.G_19_0_2\ : std_logic;
signal \Lab_UT.dictrl.nextStateZ0Z_2_cascade_\ : std_logic;
signal \Lab_UT.dictrl.dicLdASones_rst\ : std_logic;
signal \Lab_UT.dictrl.dicLdASones_rst_cascade_\ : std_logic;
signal \Lab_UT.dictrl.dicLdASonesZ0\ : std_logic;
signal \Lab_UT.dictrl.N_5ctr\ : std_logic;
signal \Lab_UT.dictrl.N_7ctr\ : std_logic;
signal \Lab_UT.dictrl.nextState_RNIGHD18Z0Z_1\ : std_logic;
signal \Lab_UT.dictrl.i8_mux\ : std_logic;
signal \Lab_UT.dictrl.currState_2_RNI1O2A_0Z0Z_1\ : std_logic;
signal \Lab_UT.dictrl.r_dicLdMtens15_1i_cascade_\ : std_logic;
signal \Lab_UT.dictrl.currState_ret_3and\ : std_logic;
signal \Lab_UT.dictrl.currState_0_ret_28_RNOZ0Z_2\ : std_logic;
signal \Lab_UT.dictrl.N_8ctr\ : std_logic;
signal \Lab_UT.dictrl.currState_0_ret_28_RNOZ0Z_3_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_8_0\ : std_logic;
signal \Lab_UT.dictrl.r_dicLdMtens21_1_reti\ : std_logic;
signal \Lab_UT.dictrl.decoder.de_littleA_2Z0Z_0\ : std_logic;
signal \Lab_UT.dictrl.de_littleA_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_37_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g0_15_rn_1\ : std_logic;
signal \Lab_UT.dictrl.G_19_0_a7_0_1\ : std_logic;
signal \G_19_0_a7_4_7\ : std_logic;
signal \Lab_UT.dictrl.currState_2_RNIEPCJZ0Z_1\ : std_logic;
signal \Lab_UT.dictrl.nextState_0_3\ : std_logic;
signal \Lab_UT.dictrl.N_1612_0\ : std_logic;
signal \Lab_UT.dictrl.currState_2_RNI2P2AZ0Z_2\ : std_logic;
signal \Lab_UT_dictrl_currState_1\ : std_logic;
signal \Lab_UT.dictrl.G_19_0_a7_2\ : std_logic;
signal \Lab_UT.dictrl.decoder.g0_2Z0Z_2\ : std_logic;
signal \Lab_UT_dictrl_decoder_de_cr_2_cascade_\ : std_logic;
signal \buart__rx_bitcount_2_rep1\ : std_logic;
signal \Lab_UT.dictrl.decoder.g0_4_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.de_cr_1_0\ : std_logic;
signal \Lab_UT.dictrl.de_cr_0\ : std_logic;
signal bu_rx_data_fast_2 : std_logic;
signal \Lab_UT.dictrl.decoder.g0_3Z0Z_0\ : std_logic;
signal \Lab_UT.dictrl.de_cr_1_2\ : std_logic;
signal \Lab_UT.dictrl.decoder.g0_4Z0Z_3\ : std_logic;
signal \Lab_UT.dictrl.decoder.g0_3_2_cascade_\ : std_logic;
signal \Lab_UT_dictrl_decoder_de_cr_1_1\ : std_logic;
signal \Lab_UT.dictrl.de_cr_2_0\ : std_logic;
signal \Lab_UT.dictrl.decoder.g0_4_1\ : std_logic;
signal \buart__rx_bitcount_4\ : std_logic;
signal \buart__rx_bitcount_3\ : std_logic;
signal \buart__rx_bitcount_2\ : std_logic;
signal \Lab_UT.dictrl.g0_8_cascade_\ : std_logic;
signal \buart__rx_valid_2_0\ : std_logic;
signal \Lab_UT.dictrl.g0_11\ : std_logic;
signal \Lab_UT.uu0.un99_ci_0_cascade_\ : std_logic;
signal \Lab_UT.uu0.un88_ci_3\ : std_logic;
signal \Lab_UT.uu0.un88_ci_3_cascade_\ : std_logic;
signal \Lab_UT.uu0.l_countZ0Z_7\ : std_logic;
signal \Lab_UT.uu0.l_countZ0Z_17\ : std_logic;
signal \Lab_UT.uu0.un110_ci_cascade_\ : std_logic;
signal \Lab_UT.uu0.un220_ci\ : std_logic;
signal \Lab_UT.uu0.l_countZ0Z_9\ : std_logic;
signal \Lab_UT.uu0.l_countZ0Z_10\ : std_logic;
signal \Lab_UT.uu0.un4_l_count_14_cascade_\ : std_logic;
signal \Lab_UT.uu0.un187_ci_1_cascade_\ : std_logic;
signal \Lab_UT.uu0.un154_ci_9\ : std_logic;
signal \Lab_UT.uu0.l_countZ0Z_14\ : std_logic;
signal \Lab_UT.uu0.un4_l_count_0_8\ : std_logic;
signal \Lab_UT.uu0.un198_ci_2\ : std_logic;
signal \Lab_UT.uu0.un110_ci\ : std_logic;
signal \Lab_UT.uu0.l_countZ0Z_8\ : std_logic;
signal \uu2.un28_w_addr_user_i_0\ : std_logic;
signal \uu2.un1_w_user_lf_0_cascade_\ : std_logic;
signal \uu2.vram_wr_en_0_iZ0\ : std_logic;
signal \uu2.un1_w_user_lf_0\ : std_logic;
signal \uu2.un3_w_addr_user\ : std_logic;
signal \uu2.un1_w_user_cr_0\ : std_logic;
signal \uu2.un1_w_user_cr_0_cascade_\ : std_logic;
signal \uu2.N_71\ : std_logic;
signal \uu2.un4_w_user_data_rdyZ0Z_0_cascade_\ : std_logic;
signal \uu2.mem0.w_data_6\ : std_logic;
signal \uu2.un1_w_user_crZ0Z_4\ : std_logic;
signal \uu2.un1_w_user_lfZ0Z_4\ : std_logic;
signal \uu2.mem0.w_data_2\ : std_logic;
signal \uu2.un4_w_user_data_rdyZ0Z_0\ : std_logic;
signal \uu2.mem0.w_addr_0\ : std_logic;
signal \INVuu2.w_addr_user_0C_net\ : std_logic;
signal \uu2.w_addr_userZ0Z_0\ : std_logic;
signal \uu2.w_addr_userZ0Z_2\ : std_logic;
signal \uu2.w_addr_userZ0Z_3\ : std_logic;
signal \uu2.w_addr_userZ0Z_1\ : std_logic;
signal \resetGen.un252_ci_cascade_\ : std_logic;
signal \resetGen.reset_countZ0Z_3\ : std_logic;
signal \resetGen.reset_countZ0Z_1\ : std_logic;
signal \resetGen.reset_countZ0Z_0\ : std_logic;
signal \resetGen.un241_ci\ : std_logic;
signal \resetGen.reset_countZ0Z_4\ : std_logic;
signal \resetGen.un241_ci_cascade_\ : std_logic;
signal \resetGen.reset_countZ0Z_2\ : std_logic;
signal \Lab_UT.uu0.delay_lineZ0Z_1\ : std_logic;
signal \Lab_UT.uu0.un11_l_count_i\ : std_logic;
signal \Lab_UT.L3_segment1_1_0_3\ : std_logic;
signal \Lab_UT.L3_segment1_0_i_1_0_cascade_\ : std_logic;
signal \uu2.bitmapZ0Z_58\ : std_logic;
signal \Lab_UT.L3_segment1_0_i_1_1\ : std_logic;
signal \Lab_UT.dictrl.enableSeg1\ : std_logic;
signal \Lab_UT.L3_segment1_1_2_cascade_\ : std_logic;
signal \INVuu2.bitmap_93C_net\ : std_logic;
signal \uu2.bitmapZ0Z_93\ : std_logic;
signal \uu2.bitmap_pmux_25_bm_1\ : std_logic;
signal \uu2.bitmapZ0Z_221\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_0\ : std_logic;
signal \uu2.bitmap_RNI1D952Z0Z_93\ : std_logic;
signal \Lab_UT.Sone_at_0\ : std_logic;
signal \Lab_UT.Sone_at_0_cascade_\ : std_logic;
signal \Lab_UT.N_77_2\ : std_logic;
signal \Lab_UT.Sone_at_3\ : std_logic;
signal \Lab_UT.Sone_at_2\ : std_logic;
signal \Lab_UT.Sten_at_1\ : std_logic;
signal \Lab_UT.Sten_at_0\ : std_logic;
signal \Lab_UT.Sten_at_3\ : std_logic;
signal \Lab_UT.Sten_at_1_cascade_\ : std_logic;
signal \Lab_UT.Sten_at_2\ : std_logic;
signal \Lab_UT.segmentUQ_0_0_0\ : std_logic;
signal \Lab_UT.dictrl.L3_segment1_1\ : std_logic;
signal \Lab_UT.Sone_at_1\ : std_logic;
signal \Lab_UT.dictrl.r_enable1_2_i_m\ : std_logic;
signal \Lab_UT.alarm_or_time_0\ : std_logic;
signal \Lab_UT.alarm_or_time_0_cascade_\ : std_logic;
signal \Lab_UT.Mten_at_2\ : std_logic;
signal \Lab_UT.dictrl.r_enable1_2_m\ : std_logic;
signal \Lab_UT.dictrl.r_enable1_2_m_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g0_i_a4_0\ : std_logic;
signal \Lab_UT.dictrl.r_enableZ0Z2\ : std_logic;
signal \Lab_UT.dictrl.enableSeg2\ : std_logic;
signal \Lab_UT.dictrl.currState_0_ret_20and_1_0\ : std_logic;
signal \Lab_UT.dictrl.r_dicLdMtens16_reti\ : std_logic;
signal \Lab_UT.dictrl.r_dicLdMtens19\ : std_logic;
signal \Lab_UT.dictrl.r_dicLdMtens22_i_6\ : std_logic;
signal \Lab_UT.dictrl.r_enable2_3_iv_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.r_enable2_3_iv_3\ : std_logic;
signal \Lab_UT.dictrl.r_Sone_init17_4\ : std_logic;
signal \Lab_UT.dictrl.r_dicLdMtens23_i_6\ : std_logic;
signal \Lab_UT.dictrl.un1_r_dicLdMtens19_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.r_alarm_or_timeZ0\ : std_logic;
signal \Lab_UT.dictrl.r_dicLdMtens18_i_6\ : std_logic;
signal \Lab_UT.dictrl.r_dicLdMtens17_i_6\ : std_logic;
signal \Lab_UT.dictrl.r_dicLdMtens16\ : std_logic;
signal \Lab_UT.dictrl.nextStateZ0Z_2\ : std_logic;
signal \Lab_UT.dictrl.nextStateZ0Z_1\ : std_logic;
signal \Lab_UT.dictrl.r_dicLdMtens17\ : std_logic;
signal \Lab_UT.dictrl.currState_ret_1and\ : std_logic;
signal \Lab_UT.dictrl.dicLdAMones_rst\ : std_logic;
signal \Lab_UT.dictrl.dicLdAMonesZ0\ : std_logic;
signal \Lab_UT.dictrl.dicLdAMones_rst_cascade_\ : std_logic;
signal \Lab_UT.dictrl.r_dicLdMtens23_2\ : std_logic;
signal \Lab_UT.dictrl.dicLdAStensZ0\ : std_logic;
signal \Lab_UT.dictrl.dicLdAStens_rst\ : std_logic;
signal \resetGen.escKeyZ0\ : std_logic;
signal \Lab_UT.dictrl.currState_3_rep1\ : std_logic;
signal \Lab_UT.dictrl.N_5\ : std_logic;
signal \Lab_UT.dictrl.N_6\ : std_logic;
signal \Lab_UT.dictrl.r_dicLdMtens14_i_6\ : std_logic;
signal \Lab_UT.dictrl.r_dicLdMtens20_i_6\ : std_logic;
signal \Lab_UT.dictrl.r_enable3_3_iv_1\ : std_logic;
signal \buart.Z_rx.G_30_0_o3_1_0_cascade_\ : std_logic;
signal \Lab_UT_dictrl_decoder_de_cr_1\ : std_logic;
signal \Lab_UT.dictrl.currStateZ0Z_0\ : std_logic;
signal \N_6_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_21_0\ : std_logic;
signal \resetGen.escKey_4_0\ : std_logic;
signal \Lab_UT.dictrl.nextStateZ0Z_0\ : std_logic;
signal \Lab_UT.dictrl.currState_0_rep2\ : std_logic;
signal \Lab_UT.dictrl.g0_7_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g0_10\ : std_logic;
signal bu_rx_data_fast_1 : std_logic;
signal bu_rx_data_3_rep1 : std_logic;
signal \Lab_UT.dictrl.g1_5_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g1_7_1\ : std_logic;
signal bu_rx_data_2_rep1 : std_logic;
signal \Lab_UT.dictrl.g1_4_1\ : std_logic;
signal \Lab_UT.dictrl.currState_fast_3\ : std_logic;
signal \buart.Z_rx.G_30_0_o3_1_4\ : std_logic;
signal \Lab_UT.dictrl.nextStateZ0Z_3\ : std_logic;
signal bu_rx_data_4_rep1 : std_logic;
signal bu_rx_data_1_rep1 : std_logic;
signal \Lab_UT.dictrl.decoder.g0Z0Z_3\ : std_logic;
signal bu_rx_data_0_rep1 : std_logic;
signal bu_rx_data_6_rep1 : std_logic;
signal bu_rx_data_5_rep1 : std_logic;
signal bu_rx_data_fast_3 : std_logic;
signal \buart.Z_rx.hhZ0Z_1\ : std_logic;
signal bu_rx_data_7_rep1 : std_logic;
signal \Lab_UT.uu0.un44_ci\ : std_logic;
signal \Lab_UT.uu0.un44_ci_cascade_\ : std_logic;
signal \Lab_UT.uu0.l_countZ0Z_3\ : std_logic;
signal \Lab_UT.uu0.l_countZ0Z_2\ : std_logic;
signal \Lab_UT.uu0.un66_ci_cascade_\ : std_logic;
signal \Lab_UT.uu0.l_countZ0Z_4\ : std_logic;
signal \Lab_UT.uu0.un66_ci\ : std_logic;
signal \Lab_UT.uu0.un11_l_count_i_g\ : std_logic;
signal \Lab_UT.uu0.delay_lineZ0Z_0\ : std_logic;
signal \Lab_UT.uu0.l_countZ0Z_5\ : std_logic;
signal \Lab_UT.uu0.l_precountZ0Z_3\ : std_logic;
signal \Lab_UT.uu0.l_countZ0Z_1\ : std_logic;
signal \Lab_UT.uu0.l_countZ0Z_18\ : std_logic;
signal \Lab_UT.uu0.l_countZ0Z_15\ : std_logic;
signal \Lab_UT.uu0.un4_l_count_11_cascade_\ : std_logic;
signal \Lab_UT.uu0.l_countZ0Z_6\ : std_logic;
signal \Lab_UT.uu0.un4_l_count_12\ : std_logic;
signal \Lab_UT.uu0.un4_l_count_16_cascade_\ : std_logic;
signal \Lab_UT.uu0.un4_l_count_18\ : std_logic;
signal \Lab_UT.uu0.l_precountZ0Z_1\ : std_logic;
signal \Lab_UT.uu0.l_countZ0Z_16\ : std_logic;
signal \Lab_UT.uu0.l_countZ0Z_11\ : std_logic;
signal \Lab_UT.uu0.l_precountZ0Z_2\ : std_logic;
signal \Lab_UT.uu0.l_countZ0Z_0\ : std_logic;
signal \Lab_UT.uu0.un4_l_count_13\ : std_logic;
signal \uu2.w_addr_userZ0Z_5\ : std_logic;
signal \uu2.w_addr_userZ0Z_4\ : std_logic;
signal \uu2.un28_w_addr_user_i\ : std_logic;
signal \uu2.un404_ci\ : std_logic;
signal \uu2.un426_ci_3\ : std_logic;
signal \uu2.w_addr_userZ0Z_6\ : std_logic;
signal \INVuu2.w_addr_user_5C_net\ : std_logic;
signal \uu2.w_addr_user_RNIMJ3O2Z0Z_2\ : std_logic;
signal \L3_tx_data_rdy\ : std_logic;
signal \L3_tx_data_6\ : std_logic;
signal \Lab_UT.display.N_88_cascade_\ : std_logic;
signal \L3_tx_data_1\ : std_logic;
signal \Lab_UT.display.N_120_cascade_\ : std_logic;
signal \L3_tx_data_4\ : std_logic;
signal \L3_tx_data_5\ : std_logic;
signal \Lab_UT.display.N_153_cascade_\ : std_logic;
signal \Lab_UT.display.dOutP_0_iv_i_1_1\ : std_logic;
signal \Lab_UT.display.N_150\ : std_logic;
signal \Lab_UT.display.N_101_cascade_\ : std_logic;
signal \Lab_UT.display.N_88\ : std_logic;
signal \Lab_UT.display.dOutP_0_iv_i_0_3_cascade_\ : std_logic;
signal \Lab_UT.display.dOutP_0_iv_i_2_3\ : std_logic;
signal \L3_tx_data_3\ : std_logic;
signal \uu2.r_addrZ0Z_5\ : std_logic;
signal \Lab_UT.di_AMones_0\ : std_logic;
signal \Lab_UT.di_AMones_2\ : std_logic;
signal \Lab_UT.ld_enable_AMones\ : std_logic;
signal \Lab_UT.di_AMones_3\ : std_logic;
signal \Lab_UT.di_ASones_0\ : std_logic;
signal \Lab_UT.di_ASones_1\ : std_logic;
signal \Lab_UT.di_ASones_2\ : std_logic;
signal \Lab_UT.ld_enable_AMtens\ : std_logic;
signal \Lab_UT.di_AStens_3\ : std_logic;
signal \Lab_UT.ld_enable_ASones\ : std_logic;
signal \Lab_UT.di_ASones_3\ : std_logic;
signal \Lab_UT.ld_enable_AStens\ : std_logic;
signal \Lab_UT.uu0.un4_l_count_0\ : std_logic;
signal \Lab_UT.halfPulse\ : std_logic;
signal \Lab_UT.displayAlarmZ0Z_1\ : std_logic;
signal \Lab_UT.dicLdStens\ : std_logic;
signal \Lab_UT.dicLdStens_latmux\ : std_logic;
signal \Lab_UT.didp.Stens_subtractor.un1_q_axb0\ : std_logic;
signal \Lab_UT.didp.Stens_subtractor.q_RNO_0_0_3\ : std_logic;
signal \Lab_UT.didp.Stens_subtractor.N_86\ : std_logic;
signal \Lab_UT.didp.Stens_subtractor.q_RNO_0_1_2\ : std_logic;
signal \Lab_UT.didp.q_RNIDDF11_3_cascade_\ : std_logic;
signal led_c_3 : std_logic;
signal \Lab_UT.didp.q_RNI1TVP_3\ : std_logic;
signal \Lab_UT.didp.q_RNIBBF11_2\ : std_logic;
signal \Lab_UT.didp.q_RNIVQVP_2\ : std_logic;
signal led_c_2 : std_logic;
signal \Lab_UT.dictrl.r_Sone_init5\ : std_logic;
signal \Lab_UT_dictrl_r_Sone_init17\ : std_logic;
signal \Lab_UT.dictrl.r_dicAlarmTrigZ0\ : std_logic;
signal \Lab_UT.displayAlarmZ0Z_5\ : std_logic;
signal \Lab_UT.dictrl.nextState_al_1\ : std_logic;
signal \Lab_UT.dictrl.nextState_al_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.un2_dicAlarmTrig_i_6\ : std_logic;
signal \Lab_UT.dictrl.nextState_al_latmux_1\ : std_logic;
signal \Lab_UT.dictrl.nextState_al_latmux_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.nextState_alZ0Z_0\ : std_logic;
signal \Lab_UT.dictrl.un2_dicAlarmTrig\ : std_logic;
signal \Lab_UT.dictrl.N_186\ : std_logic;
signal \Lab_UT.dictrl.nextState_al_0_0\ : std_logic;
signal \Lab_UT.dictrl.N_186_cascade_\ : std_logic;
signal \Lab_UT.dictrl.nextState_al_1_0_0_1\ : std_logic;
signal \Lab_UT.dictrl.currState_alZ0Z_0\ : std_logic;
signal \Lab_UT.dictrl.currState_alZ0Z_1\ : std_logic;
signal \Lab_UT.dictrl.currState_i_5_1\ : std_logic;
signal \Lab_UT.dictrl.currState_i_5_0\ : std_logic;
signal \Lab_UT.dictrl.un1_currState_8_u_ns_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.currState_ret_7_RNI03VHZ0Z1\ : std_logic;
signal \Lab_UT.dictrl.un1_currState_inv_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.currState_0_ret_1_RNIPH7FZ0Z1\ : std_logic;
signal \Lab_UT.dictrl.r_dicLdMtens14_1\ : std_logic;
signal \Lab_UT.dictrl.r_Sone_init5_1\ : std_logic;
signal \Lab_UT.dictrl.currStateZ0Z_3\ : std_logic;
signal \Lab_UT.dictrl.un1_currState_inv_1\ : std_logic;
signal \Lab_UT.dictrl.N_201_cascade_\ : std_logic;
signal \Lab_UT.dictrl.currState_2_RNIOB6H1Z0Z_2\ : std_logic;
signal \Lab_UT.dictrl.currStateZ0Z_2\ : std_logic;
signal \Lab_UT.dictrl.currState_i_5_3\ : std_logic;
signal \Lab_UT.dictrl.r_dicRun_r_1\ : std_logic;
signal \Lab_UT.dictrl.r_dicLdMtens15_1i\ : std_logic;
signal rst : std_logic;
signal \Lab_UT.dictrl.r_dicLdMtens15_1\ : std_logic;
signal \Lab_UT.dictrl.decoder.de_atSignZ0Z_4_cascade_\ : std_logic;
signal \Lab_UT.dictrl.de_atSign\ : std_logic;
signal \Lab_UT.dictrl.de_littleA_2_cascade_\ : std_logic;
signal \Lab_UT.dictrl.de_littleL\ : std_logic;
signal bu_rx_data_5 : std_logic;
signal \Lab_UT.dictrl.de_littleL_4\ : std_logic;
signal bu_rx_data_6 : std_logic;
signal \Lab_UT.dictrl.g0_4_2\ : std_logic;
signal \Lab_UT.dictrl.de_littleA_2\ : std_logic;
signal \Lab_UT.dictrl.decoder.de_littleNZ0Z_1_cascade_\ : std_logic;
signal \Lab_UT_dictrl_decoder_de_cr_2\ : std_logic;
signal \Lab_UT.n_rdy\ : std_logic;
signal \resetGen.escKeyZ0Z_3\ : std_logic;
signal \buart.Z_rx.sample_g\ : std_logic;
signal bu_rx_data_7 : std_logic;
signal bu_rx_data_4 : std_logic;
signal \Lab_UT.dictrl.decoder.de_atSignZ0Z_5\ : std_logic;
signal \Lab_UT.uu0.l_precountZ0Z_0\ : std_logic;
signal \uu2.un404_ci_0\ : std_logic;
signal \uu2.trig_rd_is_det\ : std_logic;
signal \uu2.r_addrZ0Z_4\ : std_logic;
signal \Lab_UT.di_AMtens_0\ : std_logic;
signal \Lab_UT.displayAlarmZ0Z_0\ : std_logic;
signal \Lab_UT.di_AStens_0\ : std_logic;
signal \Lab_UT.display.N_130\ : std_logic;
signal \Lab_UT.display.dOutP_0_iv_i_0_0_cascade_\ : std_logic;
signal \Lab_UT.display.dOutP_0_iv_i_1_0\ : std_logic;
signal \L3_tx_data_0\ : std_logic;
signal \Lab_UT.display.N_153\ : std_logic;
signal \Lab_UT.displayAlarmZ1Z_2\ : std_logic;
signal \Lab_UT.di_AStens_2\ : std_logic;
signal \Lab_UT.display.dOutP_0_iv_i_0_2_cascade_\ : std_logic;
signal \Lab_UT.display.dOutP_0_iv_i_1_2\ : std_logic;
signal \L3_tx_data_2\ : std_logic;
signal \Lab_UT.display.un42_dOutP_1\ : std_logic;
signal \Lab_UT.display.cnt_RNI1STE1Z0Z_1\ : std_logic;
signal \Lab_UT.display.N_151_cascade_\ : std_logic;
signal \Lab_UT.di_AMtens_3\ : std_logic;
signal \Lab_UT.display.N_124\ : std_logic;
signal rst_g : std_logic;
signal \Lab_UT.display.N_106\ : std_logic;
signal \Lab_UT.display.N_151\ : std_logic;
signal \Lab_UT.di_AMtens_2\ : std_logic;
signal \Lab_UT.display.N_115\ : std_logic;
signal \Lab_UT.di_AStens_1\ : std_logic;
signal \Lab_UT.display.N_108_cascade_\ : std_logic;
signal \Lab_UT.di_AMones_1\ : std_logic;
signal \Lab_UT.display.dOutP_0_iv_i_0_1\ : std_logic;
signal \Lab_UT.display.N_152\ : std_logic;
signal \Lab_UT.display.cntZ0Z_1\ : std_logic;
signal \Lab_UT.display.N_92\ : std_logic;
signal \Lab_UT.display.cntZ0Z_2\ : std_logic;
signal \Lab_UT.di_AMtens_1\ : std_logic;
signal \Lab_UT.display.cntZ0Z_0\ : std_logic;
signal \Lab_UT.display.N_112\ : std_logic;
signal \Lab_UT.didp.Sones_subtractor.q_RNO_0Z0Z_3_cascade_\ : std_logic;
signal \Lab_UT.didp.Sones_subtractor.q_RNO_0_0_2\ : std_logic;
signal \Lab_UT.didp.di_Sones_2\ : std_logic;
signal \Lab_UT.didp.di_Sones_3\ : std_logic;
signal \Lab_UT.didp.Sones_subtractor.un8_Mtens_ce_cascade_\ : std_logic;
signal \o_One_Sec_Pulse\ : std_logic;
signal \uu0_sec_clkD\ : std_logic;
signal \oneSecStrb\ : std_logic;
signal \Lab_UT.ld_enable_dicRun\ : std_logic;
signal \Lab_UT.didp.N_84_cascade_\ : std_logic;
signal \Lab_UT.didp.Sones_subtractor.un8_Mtens_ce\ : std_logic;
signal \Lab_UT.didp.Stens_subtractor.q_RNI775L5_0Z0Z_3\ : std_logic;
signal \Lab_UT.didp.Stens_subtractor.q_RNI775L5_0Z0Z_3_cascade_\ : std_logic;
signal \Lab_UT.didp.Stens_subtractor.un1_q_c2\ : std_logic;
signal \Lab_UT.didp.Stens_subtractor.q_RNI8PD76Z0Z_1\ : std_logic;
signal \Lab_UT.ld_enable_Stens\ : std_logic;
signal \Lab_UT.didp.Stens_subtractor.q_7_i_1_1\ : std_logic;
signal \Lab_UT.didp.Mtens_subtractor.q_RNO_0_3_2_cascade_\ : std_logic;
signal \Lab_UT.didp.N_83\ : std_logic;
signal \Lab_UT.didp.un3_Mtens_rst_cascade_\ : std_logic;
signal \Lab_UT.didp.q_RNI775L5_3\ : std_logic;
signal \Lab_UT.didp.Mtens_subtractor.un1_q_axb0_cascade_\ : std_logic;
signal \Lab_UT.didp.Mtens_ce\ : std_logic;
signal \Lab_UT.di_Mtens_2\ : std_logic;
signal \Lab_UT.didp.Mtens_ce_cascade_\ : std_logic;
signal \Lab_UT.didp.Mtens_subtractor.q_RNO_0_2_3_cascade_\ : std_logic;
signal \Lab_UT.didp.di_Mtens_3\ : std_logic;
signal \Lab_UT.dicLdMones\ : std_logic;
signal \Lab_UT.dictrl.r_dicLdMtens14\ : std_logic;
signal \Lab_UT.dictrl.de_num0to5_1\ : std_logic;
signal \Lab_UT.dicLdMtens_latmux_cascade_\ : std_logic;
signal \Lab_UT.didp.di_Stens_2\ : std_logic;
signal \Lab_UT.didp.di_Stens_3\ : std_logic;
signal \Lab_UT.didp.un6_Mtens_ce\ : std_logic;
signal \Lab_UT.didp.un3_Mtens_rst\ : std_logic;
signal \Lab_UT.didp.Mtens_subtractor.q_RNO_2Z0Z_1\ : std_logic;
signal \Lab_UT.dicLdMtens\ : std_logic;
signal \Lab_UT.dicLdMtens_latmux\ : std_logic;
signal \Lab_UT.didp.Mtens_subtractor.N_147\ : std_logic;
signal \Lab_UT.didp.Mtens_subtractor.N_87\ : std_logic;
signal \Lab_UT.didp.Mtens_subtractor.N_145\ : std_logic;
signal \Lab_UT.didp.Mtens_subtractor.un1_q_c2\ : std_logic;
signal \Lab_UT.didp.di_Mtens_1\ : std_logic;
signal \Lab_UT.didp.q_RNITOVP_1_cascade_\ : std_logic;
signal led_c_1 : std_logic;
signal \Lab_UT.didp.di_Stens_1\ : std_logic;
signal \Lab_UT.didp.q_RNI99F11_1\ : std_logic;
signal \Lab_UT.dictrl.r_dicLdMtens15\ : std_logic;
signal bu_rx_data_rdy : std_logic;
signal \Lab_UT.dictrl.de_num_0\ : std_logic;
signal \Lab_UT.dicLdMones_latmux\ : std_logic;
signal \Lab_UT.displayAlarmZ0Z_6\ : std_logic;
signal \Lab_UT.alarm_armed\ : std_logic;
signal \Lab_UT.displayAlarmZ0Z_4\ : std_logic;
signal \Lab_UT.alarm_match\ : std_logic;
signal \Lab_UT.ld_enable_Sones_cascade_\ : std_logic;
signal \Lab_UT.didp.Sones_subtractor.q_RNO_1Z0Z_1\ : std_logic;
signal \Lab_UT.didp.Sones_subtractor.q_7_i_1_1_cascade_\ : std_logic;
signal \Lab_UT.didp.Sones_subtractor.q_RNI775L5_1_3\ : std_logic;
signal \Lab_UT.didp.N_82\ : std_logic;
signal \Lab_UT.didp.Sones_subtractor.un1_q_axb0_cascade_\ : std_logic;
signal \Lab_UT.didp.Sones_subtractor.N_85\ : std_logic;
signal \Lab_UT.didp.di_Sones_1\ : std_logic;
signal \Lab_UT.didp.N_81\ : std_logic;
signal \Lab_UT.didp.Sones_subtractor.un1_q_c2\ : std_logic;
signal \Lab_UT.didp.un4_Mtens_ce\ : std_logic;
signal \Lab_UT.didp.Mones_subtractor.un1_q_axb_0_cascade_\ : std_logic;
signal bu_rx_data_0 : std_logic;
signal bu_rx_data_3 : std_logic;
signal bu_rx_data_1 : std_logic;
signal \Lab_UT.didp.N_84\ : std_logic;
signal \Lab_UT.didp.Mones_subtractor.q_0_sqmuxa\ : std_logic;
signal \Lab_UT.didp.Mones_subtractor.q_RNO_0_2_2_cascade_\ : std_logic;
signal bu_rx_data_2 : std_logic;
signal \Lab_UT.didp.q20_0_i\ : std_logic;
signal \bfn_12_9_0_\ : std_logic;
signal \Lab_UT.didp.Mones_subtractor.un1_q_cry_0_s1\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \Lab_UT.didp.di_Mones_2\ : std_logic;
signal \Lab_UT.didp.Mones_subtractor.un1_q_cry_1_s1_THRU_CO\ : std_logic;
signal \Lab_UT.didp.Mones_subtractor.un1_q_cry_1_s1\ : std_logic;
signal \Lab_UT.didp.di_Mones_3\ : std_logic;
signal \Lab_UT.didp.Mones_subtractor.un1_q_cry_2_s1\ : std_logic;
signal \Lab_UT.didp.Mones_subtractor.q_RNO_0_1_3\ : std_logic;
signal \Lab_UT.didp.Mones_subtractor.un1_q_cry_0_s1_THRU_CO\ : std_logic;
signal \Lab_UT.didp.Mones_subtractor.N_80\ : std_logic;
signal \Lab_UT.didp.di_Mones_1\ : std_logic;
signal \Lab_UT.didp.Mones_subtractor.q_RNO_0Z0Z_1\ : std_logic;
signal \Lab_UT.didp.di_MtensZ0Z_0\ : std_logic;
signal \Lab_UT.didp.di_Mones_0\ : std_logic;
signal \Lab_UT.un1_r_Sone_init5_1_0\ : std_logic;
signal \Lab_UT.dictrl.N_258_i\ : std_logic;
signal \Lab_UT.dicLdSones_latmux\ : std_logic;
signal \Lab_UT.dicLdSones\ : std_logic;
signal \Lab_UT.didp.di_Sones_0\ : std_logic;
signal \Lab_UT.didp.curr_LEDZ0Z_0\ : std_logic;
signal \Lab_UT.didp.di_Stens_0\ : std_logic;
signal \Lab_UT.didp.q_RNIRMVP_0\ : std_logic;
signal \Lab_UT.didp.q_RNI77F11_0_cascade_\ : std_logic;
signal \Lab_UT.didp.curr_LEDZ0Z_1\ : std_logic;
signal led_c_0 : std_logic;
signal \Lab_UT.dictrl.un1_nextState_al24_0\ : std_logic;
signal \Lab_UT.alarm_off\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal clk_g : std_logic;
signal \Lab_UT.dictrl.nextState_al22\ : std_logic;

signal led_wire : std_logic_vector(4 downto 0);
signal from_pc_wire : std_logic;
signal clk_in_wire : std_logic;
signal to_ir_wire : std_logic;
signal o_serial_data_wire : std_logic;
signal sd_wire : std_logic;
signal \latticehx1k_pll_inst.latticehx1k_pll_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    led <= led_wire;
    from_pc_wire <= from_pc;
    clk_in_wire <= clk_in;
    to_ir <= to_ir_wire;
    o_serial_data <= o_serial_data_wire;
    sd <= sd_wire;
    \latticehx1k_pll_inst.latticehx1k_pll_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;
    \uu2.r_data_wire_7\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(14);
    \uu2.r_data_wire_6\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(12);
    \uu2.r_data_wire_5\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(10);
    \uu2.r_data_wire_4\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(8);
    \uu2.r_data_wire_3\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(6);
    \uu2.r_data_wire_2\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(4);
    \uu2.r_data_wire_1\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(2);
    \uu2.r_data_wire_0\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(0);
    \uu2.mem0.ram512X8_inst_physical_RADDR_wire\ <= '0'&'0'&\N__13390\&\N__13363\&\N__13696\&\N__22806\&\N__25114\&\N__13561\&\N__13669\&\N__13636\&\N__13603\;
    \uu2.mem0.ram512X8_inst_physical_WADDR_wire\ <= '0'&'0'&\N__12634\&\N__12700\&\N__14524\&\N__14536\&\N__14551\&\N__16192\&\N__14563\&\N__12685\&\N__18715\;
    \uu2.mem0.ram512X8_inst_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \uu2.mem0.ram512X8_inst_physical_WDATA_wire\ <= '0'&'0'&'0'&\N__18844\&'0'&\N__12574\&'0'&\N__12580\&'0'&\N__12559\&'0'&\N__18817\&'0'&\N__12553\&'0'&\N__12655\;

    \latticehx1k_pll_inst.latticehx1k_pll_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "110",
            DIVF => "0111111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => \latticehx1k_pll_inst.clk\,
            REFERENCECLK => \N__10939\,
            RESETB => \N__28354\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \latticehx1k_pll_inst.latticehx1k_pll_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => OPEN
        );

    \uu2.mem0.ram512X8_inst_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_F => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_E => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_D => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_C => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_B => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_A => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_9 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_8 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_7 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_6 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_5 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_4 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_3 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_2 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_1 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000"
        )
    port map (
            RDATA => \uu2.mem0.ram512X8_inst_physical_RDATA_wire\,
            RADDR => \uu2.mem0.ram512X8_inst_physical_RADDR_wire\,
            WADDR => \uu2.mem0.ram512X8_inst_physical_WADDR_wire\,
            MASK => \uu2.mem0.ram512X8_inst_physical_MASK_wire\,
            WDATA => \uu2.mem0.ram512X8_inst_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__29462\,
            RE => \N__28355\,
            WCLKE => \N__18919\,
            WCLK => \N__29461\,
            WE => \N__18918\
        );

    \led_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__30236\,
            DIN => \N__30235\,
            DOUT => \N__30234\,
            PACKAGEPIN => led_wire(1)
        );

    \led_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__30236\,
            PADOUT => \N__30235\,
            PADIN => \N__30234\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__27889\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__30227\,
            DIN => \N__30226\,
            DOUT => \N__30225\,
            PACKAGEPIN => led_wire(3)
        );

    \led_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__30227\,
            PADOUT => \N__30226\,
            PADIN => \N__30225\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__23530\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__30218\,
            DIN => \N__30217\,
            DOUT => \N__30216\,
            PACKAGEPIN => led_wire(0)
        );

    \led_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__30218\,
            PADOUT => \N__30217\,
            PADIN => \N__30216\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__29596\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \Z_rcxd.Z_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__30209\,
            DIN => \N__30208\,
            DOUT => \N__30207\,
            PACKAGEPIN => from_pc_wire
        );

    \Z_rcxd.Z_io_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000000",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__30209\,
            PADOUT => \N__30208\,
            PADIN => \N__30207\,
            CLOCKENABLE => 'H',
            DOUT1 => \GNDG0\,
            OUTPUTENABLE => '0',
            DIN0 => \uart_RXD\,
            DOUT0 => \GNDG0\,
            INPUTCLK => \N__29419\,
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \clk_in_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__30200\,
            DIN => \N__30199\,
            DOUT => \N__30198\,
            PACKAGEPIN => clk_in_wire
        );

    \clk_in_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__30200\,
            PADOUT => \N__30199\,
            PADIN => \N__30198\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => clk_in_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \to_ir_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__30191\,
            DIN => \N__30190\,
            DOUT => \N__30189\,
            PACKAGEPIN => to_ir_wire
        );

    \to_ir_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__30191\,
            PADOUT => \N__30190\,
            PADIN => \N__30189\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_serial_data_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__30182\,
            DIN => \N__30181\,
            DOUT => \N__30180\,
            PACKAGEPIN => o_serial_data_wire
        );

    \o_serial_data_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__30182\,
            PADOUT => \N__30181\,
            PADIN => \N__30180\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11923\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \sd_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__30173\,
            DIN => \N__30172\,
            DOUT => \N__30171\,
            PACKAGEPIN => sd_wire
        );

    \sd_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__30173\,
            PADOUT => \N__30172\,
            PADIN => \N__30171\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__30164\,
            DIN => \N__30163\,
            DOUT => \N__30162\,
            PACKAGEPIN => led_wire(2)
        );

    \led_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__30164\,
            PADOUT => \N__30163\,
            PADIN => \N__30162\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__23494\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__30155\,
            DIN => \N__30154\,
            DOUT => \N__30153\,
            PACKAGEPIN => led_wire(4)
        );

    \led_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__30155\,
            PADOUT => \N__30154\,
            PADIN => \N__30153\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__7323\ : CascadeMux
    port map (
            O => \N__30136\,
            I => \N__30133\
        );

    \I__7322\ : InMux
    port map (
            O => \N__30133\,
            I => \N__30130\
        );

    \I__7321\ : LocalMux
    port map (
            O => \N__30130\,
            I => \Lab_UT.didp.Mones_subtractor.q_RNO_0_1_3\
        );

    \I__7320\ : InMux
    port map (
            O => \N__30127\,
            I => \N__30124\
        );

    \I__7319\ : LocalMux
    port map (
            O => \N__30124\,
            I => \Lab_UT.didp.Mones_subtractor.un1_q_cry_0_s1_THRU_CO\
        );

    \I__7318\ : InMux
    port map (
            O => \N__30121\,
            I => \N__30113\
        );

    \I__7317\ : InMux
    port map (
            O => \N__30120\,
            I => \N__30113\
        );

    \I__7316\ : InMux
    port map (
            O => \N__30119\,
            I => \N__30108\
        );

    \I__7315\ : InMux
    port map (
            O => \N__30118\,
            I => \N__30108\
        );

    \I__7314\ : LocalMux
    port map (
            O => \N__30113\,
            I => \N__30104\
        );

    \I__7313\ : LocalMux
    port map (
            O => \N__30108\,
            I => \N__30101\
        );

    \I__7312\ : InMux
    port map (
            O => \N__30107\,
            I => \N__30098\
        );

    \I__7311\ : Span4Mux_v
    port map (
            O => \N__30104\,
            I => \N__30095\
        );

    \I__7310\ : Span4Mux_s1_h
    port map (
            O => \N__30101\,
            I => \N__30092\
        );

    \I__7309\ : LocalMux
    port map (
            O => \N__30098\,
            I => \N__30089\
        );

    \I__7308\ : Odrv4
    port map (
            O => \N__30095\,
            I => \Lab_UT.didp.Mones_subtractor.N_80\
        );

    \I__7307\ : Odrv4
    port map (
            O => \N__30092\,
            I => \Lab_UT.didp.Mones_subtractor.N_80\
        );

    \I__7306\ : Odrv12
    port map (
            O => \N__30089\,
            I => \Lab_UT.didp.Mones_subtractor.N_80\
        );

    \I__7305\ : InMux
    port map (
            O => \N__30082\,
            I => \N__30078\
        );

    \I__7304\ : InMux
    port map (
            O => \N__30081\,
            I => \N__30075\
        );

    \I__7303\ : LocalMux
    port map (
            O => \N__30078\,
            I => \N__30069\
        );

    \I__7302\ : LocalMux
    port map (
            O => \N__30075\,
            I => \N__30066\
        );

    \I__7301\ : InMux
    port map (
            O => \N__30074\,
            I => \N__30061\
        );

    \I__7300\ : InMux
    port map (
            O => \N__30073\,
            I => \N__30061\
        );

    \I__7299\ : InMux
    port map (
            O => \N__30072\,
            I => \N__30058\
        );

    \I__7298\ : Span4Mux_h
    port map (
            O => \N__30069\,
            I => \N__30055\
        );

    \I__7297\ : Odrv4
    port map (
            O => \N__30066\,
            I => \Lab_UT.didp.di_Mones_1\
        );

    \I__7296\ : LocalMux
    port map (
            O => \N__30061\,
            I => \Lab_UT.didp.di_Mones_1\
        );

    \I__7295\ : LocalMux
    port map (
            O => \N__30058\,
            I => \Lab_UT.didp.di_Mones_1\
        );

    \I__7294\ : Odrv4
    port map (
            O => \N__30055\,
            I => \Lab_UT.didp.di_Mones_1\
        );

    \I__7293\ : InMux
    port map (
            O => \N__30046\,
            I => \N__30043\
        );

    \I__7292\ : LocalMux
    port map (
            O => \N__30043\,
            I => \Lab_UT.didp.Mones_subtractor.q_RNO_0Z0Z_1\
        );

    \I__7291\ : InMux
    port map (
            O => \N__30040\,
            I => \N__30034\
        );

    \I__7290\ : InMux
    port map (
            O => \N__30039\,
            I => \N__30031\
        );

    \I__7289\ : InMux
    port map (
            O => \N__30038\,
            I => \N__30024\
        );

    \I__7288\ : InMux
    port map (
            O => \N__30037\,
            I => \N__30021\
        );

    \I__7287\ : LocalMux
    port map (
            O => \N__30034\,
            I => \N__30016\
        );

    \I__7286\ : LocalMux
    port map (
            O => \N__30031\,
            I => \N__30016\
        );

    \I__7285\ : InMux
    port map (
            O => \N__30030\,
            I => \N__30013\
        );

    \I__7284\ : InMux
    port map (
            O => \N__30029\,
            I => \N__30006\
        );

    \I__7283\ : InMux
    port map (
            O => \N__30028\,
            I => \N__30006\
        );

    \I__7282\ : InMux
    port map (
            O => \N__30027\,
            I => \N__30006\
        );

    \I__7281\ : LocalMux
    port map (
            O => \N__30024\,
            I => \N__30003\
        );

    \I__7280\ : LocalMux
    port map (
            O => \N__30021\,
            I => \Lab_UT.didp.di_MtensZ0Z_0\
        );

    \I__7279\ : Odrv4
    port map (
            O => \N__30016\,
            I => \Lab_UT.didp.di_MtensZ0Z_0\
        );

    \I__7278\ : LocalMux
    port map (
            O => \N__30013\,
            I => \Lab_UT.didp.di_MtensZ0Z_0\
        );

    \I__7277\ : LocalMux
    port map (
            O => \N__30006\,
            I => \Lab_UT.didp.di_MtensZ0Z_0\
        );

    \I__7276\ : Odrv12
    port map (
            O => \N__30003\,
            I => \Lab_UT.didp.di_MtensZ0Z_0\
        );

    \I__7275\ : InMux
    port map (
            O => \N__29992\,
            I => \N__29989\
        );

    \I__7274\ : LocalMux
    port map (
            O => \N__29989\,
            I => \N__29982\
        );

    \I__7273\ : InMux
    port map (
            O => \N__29988\,
            I => \N__29977\
        );

    \I__7272\ : InMux
    port map (
            O => \N__29987\,
            I => \N__29977\
        );

    \I__7271\ : InMux
    port map (
            O => \N__29986\,
            I => \N__29972\
        );

    \I__7270\ : InMux
    port map (
            O => \N__29985\,
            I => \N__29972\
        );

    \I__7269\ : Span4Mux_h
    port map (
            O => \N__29982\,
            I => \N__29969\
        );

    \I__7268\ : LocalMux
    port map (
            O => \N__29977\,
            I => \Lab_UT.didp.di_Mones_0\
        );

    \I__7267\ : LocalMux
    port map (
            O => \N__29972\,
            I => \Lab_UT.didp.di_Mones_0\
        );

    \I__7266\ : Odrv4
    port map (
            O => \N__29969\,
            I => \Lab_UT.didp.di_Mones_0\
        );

    \I__7265\ : CascadeMux
    port map (
            O => \N__29962\,
            I => \N__29953\
        );

    \I__7264\ : InMux
    port map (
            O => \N__29961\,
            I => \N__29945\
        );

    \I__7263\ : InMux
    port map (
            O => \N__29960\,
            I => \N__29945\
        );

    \I__7262\ : InMux
    port map (
            O => \N__29959\,
            I => \N__29940\
        );

    \I__7261\ : InMux
    port map (
            O => \N__29958\,
            I => \N__29940\
        );

    \I__7260\ : InMux
    port map (
            O => \N__29957\,
            I => \N__29936\
        );

    \I__7259\ : InMux
    port map (
            O => \N__29956\,
            I => \N__29929\
        );

    \I__7258\ : InMux
    port map (
            O => \N__29953\,
            I => \N__29929\
        );

    \I__7257\ : InMux
    port map (
            O => \N__29952\,
            I => \N__29929\
        );

    \I__7256\ : InMux
    port map (
            O => \N__29951\,
            I => \N__29924\
        );

    \I__7255\ : InMux
    port map (
            O => \N__29950\,
            I => \N__29924\
        );

    \I__7254\ : LocalMux
    port map (
            O => \N__29945\,
            I => \N__29921\
        );

    \I__7253\ : LocalMux
    port map (
            O => \N__29940\,
            I => \N__29918\
        );

    \I__7252\ : InMux
    port map (
            O => \N__29939\,
            I => \N__29915\
        );

    \I__7251\ : LocalMux
    port map (
            O => \N__29936\,
            I => \N__29912\
        );

    \I__7250\ : LocalMux
    port map (
            O => \N__29929\,
            I => \N__29905\
        );

    \I__7249\ : LocalMux
    port map (
            O => \N__29924\,
            I => \N__29905\
        );

    \I__7248\ : Span4Mux_v
    port map (
            O => \N__29921\,
            I => \N__29905\
        );

    \I__7247\ : Span4Mux_s3_h
    port map (
            O => \N__29918\,
            I => \N__29902\
        );

    \I__7246\ : LocalMux
    port map (
            O => \N__29915\,
            I => \Lab_UT.un1_r_Sone_init5_1_0\
        );

    \I__7245\ : Odrv12
    port map (
            O => \N__29912\,
            I => \Lab_UT.un1_r_Sone_init5_1_0\
        );

    \I__7244\ : Odrv4
    port map (
            O => \N__29905\,
            I => \Lab_UT.un1_r_Sone_init5_1_0\
        );

    \I__7243\ : Odrv4
    port map (
            O => \N__29902\,
            I => \Lab_UT.un1_r_Sone_init5_1_0\
        );

    \I__7242\ : InMux
    port map (
            O => \N__29893\,
            I => \N__29888\
        );

    \I__7241\ : InMux
    port map (
            O => \N__29892\,
            I => \N__29883\
        );

    \I__7240\ : InMux
    port map (
            O => \N__29891\,
            I => \N__29883\
        );

    \I__7239\ : LocalMux
    port map (
            O => \N__29888\,
            I => \N__29877\
        );

    \I__7238\ : LocalMux
    port map (
            O => \N__29883\,
            I => \N__29877\
        );

    \I__7237\ : InMux
    port map (
            O => \N__29882\,
            I => \N__29874\
        );

    \I__7236\ : Odrv12
    port map (
            O => \N__29877\,
            I => \Lab_UT.dictrl.N_258_i\
        );

    \I__7235\ : LocalMux
    port map (
            O => \N__29874\,
            I => \Lab_UT.dictrl.N_258_i\
        );

    \I__7234\ : InMux
    port map (
            O => \N__29869\,
            I => \N__29864\
        );

    \I__7233\ : InMux
    port map (
            O => \N__29868\,
            I => \N__29859\
        );

    \I__7232\ : InMux
    port map (
            O => \N__29867\,
            I => \N__29859\
        );

    \I__7231\ : LocalMux
    port map (
            O => \N__29864\,
            I => \N__29854\
        );

    \I__7230\ : LocalMux
    port map (
            O => \N__29859\,
            I => \N__29854\
        );

    \I__7229\ : Span4Mux_v
    port map (
            O => \N__29854\,
            I => \N__29851\
        );

    \I__7228\ : Span4Mux_h
    port map (
            O => \N__29851\,
            I => \N__29848\
        );

    \I__7227\ : Odrv4
    port map (
            O => \N__29848\,
            I => \Lab_UT.dicLdSones_latmux\
        );

    \I__7226\ : CascadeMux
    port map (
            O => \N__29845\,
            I => \N__29840\
        );

    \I__7225\ : CascadeMux
    port map (
            O => \N__29844\,
            I => \N__29837\
        );

    \I__7224\ : InMux
    port map (
            O => \N__29843\,
            I => \N__29832\
        );

    \I__7223\ : InMux
    port map (
            O => \N__29840\,
            I => \N__29832\
        );

    \I__7222\ : InMux
    port map (
            O => \N__29837\,
            I => \N__29829\
        );

    \I__7221\ : LocalMux
    port map (
            O => \N__29832\,
            I => \N__29826\
        );

    \I__7220\ : LocalMux
    port map (
            O => \N__29829\,
            I => \Lab_UT.dicLdSones\
        );

    \I__7219\ : Odrv12
    port map (
            O => \N__29826\,
            I => \Lab_UT.dicLdSones\
        );

    \I__7218\ : InMux
    port map (
            O => \N__29821\,
            I => \N__29817\
        );

    \I__7217\ : InMux
    port map (
            O => \N__29820\,
            I => \N__29809\
        );

    \I__7216\ : LocalMux
    port map (
            O => \N__29817\,
            I => \N__29806\
        );

    \I__7215\ : InMux
    port map (
            O => \N__29816\,
            I => \N__29799\
        );

    \I__7214\ : InMux
    port map (
            O => \N__29815\,
            I => \N__29799\
        );

    \I__7213\ : InMux
    port map (
            O => \N__29814\,
            I => \N__29799\
        );

    \I__7212\ : InMux
    port map (
            O => \N__29813\,
            I => \N__29794\
        );

    \I__7211\ : InMux
    port map (
            O => \N__29812\,
            I => \N__29794\
        );

    \I__7210\ : LocalMux
    port map (
            O => \N__29809\,
            I => \N__29791\
        );

    \I__7209\ : Odrv4
    port map (
            O => \N__29806\,
            I => \Lab_UT.didp.di_Sones_0\
        );

    \I__7208\ : LocalMux
    port map (
            O => \N__29799\,
            I => \Lab_UT.didp.di_Sones_0\
        );

    \I__7207\ : LocalMux
    port map (
            O => \N__29794\,
            I => \Lab_UT.didp.di_Sones_0\
        );

    \I__7206\ : Odrv12
    port map (
            O => \N__29791\,
            I => \Lab_UT.didp.di_Sones_0\
        );

    \I__7205\ : InMux
    port map (
            O => \N__29782\,
            I => \N__29775\
        );

    \I__7204\ : InMux
    port map (
            O => \N__29781\,
            I => \N__29768\
        );

    \I__7203\ : InMux
    port map (
            O => \N__29780\,
            I => \N__29768\
        );

    \I__7202\ : CascadeMux
    port map (
            O => \N__29779\,
            I => \N__29765\
        );

    \I__7201\ : CascadeMux
    port map (
            O => \N__29778\,
            I => \N__29762\
        );

    \I__7200\ : LocalMux
    port map (
            O => \N__29775\,
            I => \N__29758\
        );

    \I__7199\ : InMux
    port map (
            O => \N__29774\,
            I => \N__29755\
        );

    \I__7198\ : InMux
    port map (
            O => \N__29773\,
            I => \N__29752\
        );

    \I__7197\ : LocalMux
    port map (
            O => \N__29768\,
            I => \N__29749\
        );

    \I__7196\ : InMux
    port map (
            O => \N__29765\,
            I => \N__29744\
        );

    \I__7195\ : InMux
    port map (
            O => \N__29762\,
            I => \N__29744\
        );

    \I__7194\ : InMux
    port map (
            O => \N__29761\,
            I => \N__29741\
        );

    \I__7193\ : Span4Mux_v
    port map (
            O => \N__29758\,
            I => \N__29736\
        );

    \I__7192\ : LocalMux
    port map (
            O => \N__29755\,
            I => \N__29736\
        );

    \I__7191\ : LocalMux
    port map (
            O => \N__29752\,
            I => \N__29733\
        );

    \I__7190\ : Span4Mux_s3_h
    port map (
            O => \N__29749\,
            I => \N__29726\
        );

    \I__7189\ : LocalMux
    port map (
            O => \N__29744\,
            I => \N__29726\
        );

    \I__7188\ : LocalMux
    port map (
            O => \N__29741\,
            I => \N__29726\
        );

    \I__7187\ : Span4Mux_v
    port map (
            O => \N__29736\,
            I => \N__29721\
        );

    \I__7186\ : Span4Mux_v
    port map (
            O => \N__29733\,
            I => \N__29718\
        );

    \I__7185\ : Span4Mux_v
    port map (
            O => \N__29726\,
            I => \N__29715\
        );

    \I__7184\ : InMux
    port map (
            O => \N__29725\,
            I => \N__29710\
        );

    \I__7183\ : InMux
    port map (
            O => \N__29724\,
            I => \N__29710\
        );

    \I__7182\ : Odrv4
    port map (
            O => \N__29721\,
            I => \Lab_UT.didp.curr_LEDZ0Z_0\
        );

    \I__7181\ : Odrv4
    port map (
            O => \N__29718\,
            I => \Lab_UT.didp.curr_LEDZ0Z_0\
        );

    \I__7180\ : Odrv4
    port map (
            O => \N__29715\,
            I => \Lab_UT.didp.curr_LEDZ0Z_0\
        );

    \I__7179\ : LocalMux
    port map (
            O => \N__29710\,
            I => \Lab_UT.didp.curr_LEDZ0Z_0\
        );

    \I__7178\ : InMux
    port map (
            O => \N__29701\,
            I => \N__29696\
        );

    \I__7177\ : InMux
    port map (
            O => \N__29700\,
            I => \N__29693\
        );

    \I__7176\ : InMux
    port map (
            O => \N__29699\,
            I => \N__29690\
        );

    \I__7175\ : LocalMux
    port map (
            O => \N__29696\,
            I => \N__29686\
        );

    \I__7174\ : LocalMux
    port map (
            O => \N__29693\,
            I => \N__29678\
        );

    \I__7173\ : LocalMux
    port map (
            O => \N__29690\,
            I => \N__29678\
        );

    \I__7172\ : InMux
    port map (
            O => \N__29689\,
            I => \N__29675\
        );

    \I__7171\ : Span4Mux_v
    port map (
            O => \N__29686\,
            I => \N__29672\
        );

    \I__7170\ : InMux
    port map (
            O => \N__29685\,
            I => \N__29665\
        );

    \I__7169\ : InMux
    port map (
            O => \N__29684\,
            I => \N__29665\
        );

    \I__7168\ : InMux
    port map (
            O => \N__29683\,
            I => \N__29665\
        );

    \I__7167\ : Span4Mux_s3_h
    port map (
            O => \N__29678\,
            I => \N__29660\
        );

    \I__7166\ : LocalMux
    port map (
            O => \N__29675\,
            I => \N__29660\
        );

    \I__7165\ : Odrv4
    port map (
            O => \N__29672\,
            I => \Lab_UT.didp.di_Stens_0\
        );

    \I__7164\ : LocalMux
    port map (
            O => \N__29665\,
            I => \Lab_UT.didp.di_Stens_0\
        );

    \I__7163\ : Odrv4
    port map (
            O => \N__29660\,
            I => \Lab_UT.didp.di_Stens_0\
        );

    \I__7162\ : InMux
    port map (
            O => \N__29653\,
            I => \N__29650\
        );

    \I__7161\ : LocalMux
    port map (
            O => \N__29650\,
            I => \Lab_UT.didp.q_RNIRMVP_0\
        );

    \I__7160\ : CascadeMux
    port map (
            O => \N__29647\,
            I => \Lab_UT.didp.q_RNI77F11_0_cascade_\
        );

    \I__7159\ : InMux
    port map (
            O => \N__29644\,
            I => \N__29641\
        );

    \I__7158\ : LocalMux
    port map (
            O => \N__29641\,
            I => \N__29638\
        );

    \I__7157\ : Span4Mux_v
    port map (
            O => \N__29638\,
            I => \N__29634\
        );

    \I__7156\ : InMux
    port map (
            O => \N__29637\,
            I => \N__29631\
        );

    \I__7155\ : IoSpan4Mux
    port map (
            O => \N__29634\,
            I => \N__29624\
        );

    \I__7154\ : LocalMux
    port map (
            O => \N__29631\,
            I => \N__29624\
        );

    \I__7153\ : InMux
    port map (
            O => \N__29630\,
            I => \N__29619\
        );

    \I__7152\ : InMux
    port map (
            O => \N__29629\,
            I => \N__29619\
        );

    \I__7151\ : Span4Mux_s3_h
    port map (
            O => \N__29624\,
            I => \N__29616\
        );

    \I__7150\ : LocalMux
    port map (
            O => \N__29619\,
            I => \N__29613\
        );

    \I__7149\ : Span4Mux_v
    port map (
            O => \N__29616\,
            I => \N__29609\
        );

    \I__7148\ : Span4Mux_v
    port map (
            O => \N__29613\,
            I => \N__29606\
        );

    \I__7147\ : InMux
    port map (
            O => \N__29612\,
            I => \N__29603\
        );

    \I__7146\ : Odrv4
    port map (
            O => \N__29609\,
            I => \Lab_UT.didp.curr_LEDZ0Z_1\
        );

    \I__7145\ : Odrv4
    port map (
            O => \N__29606\,
            I => \Lab_UT.didp.curr_LEDZ0Z_1\
        );

    \I__7144\ : LocalMux
    port map (
            O => \N__29603\,
            I => \Lab_UT.didp.curr_LEDZ0Z_1\
        );

    \I__7143\ : IoInMux
    port map (
            O => \N__29596\,
            I => \N__29593\
        );

    \I__7142\ : LocalMux
    port map (
            O => \N__29593\,
            I => \N__29590\
        );

    \I__7141\ : Span4Mux_s0_h
    port map (
            O => \N__29590\,
            I => \N__29587\
        );

    \I__7140\ : Odrv4
    port map (
            O => \N__29587\,
            I => led_c_0
        );

    \I__7139\ : InMux
    port map (
            O => \N__29584\,
            I => \N__29581\
        );

    \I__7138\ : LocalMux
    port map (
            O => \N__29581\,
            I => \N__29578\
        );

    \I__7137\ : Span4Mux_s2_h
    port map (
            O => \N__29578\,
            I => \N__29569\
        );

    \I__7136\ : InMux
    port map (
            O => \N__29577\,
            I => \N__29562\
        );

    \I__7135\ : InMux
    port map (
            O => \N__29576\,
            I => \N__29562\
        );

    \I__7134\ : InMux
    port map (
            O => \N__29575\,
            I => \N__29562\
        );

    \I__7133\ : InMux
    port map (
            O => \N__29574\,
            I => \N__29555\
        );

    \I__7132\ : InMux
    port map (
            O => \N__29573\,
            I => \N__29555\
        );

    \I__7131\ : InMux
    port map (
            O => \N__29572\,
            I => \N__29555\
        );

    \I__7130\ : Odrv4
    port map (
            O => \N__29569\,
            I => \Lab_UT.dictrl.un1_nextState_al24_0\
        );

    \I__7129\ : LocalMux
    port map (
            O => \N__29562\,
            I => \Lab_UT.dictrl.un1_nextState_al24_0\
        );

    \I__7128\ : LocalMux
    port map (
            O => \N__29555\,
            I => \Lab_UT.dictrl.un1_nextState_al24_0\
        );

    \I__7127\ : InMux
    port map (
            O => \N__29548\,
            I => \N__29541\
        );

    \I__7126\ : InMux
    port map (
            O => \N__29547\,
            I => \N__29541\
        );

    \I__7125\ : InMux
    port map (
            O => \N__29546\,
            I => \N__29536\
        );

    \I__7124\ : LocalMux
    port map (
            O => \N__29541\,
            I => \N__29533\
        );

    \I__7123\ : InMux
    port map (
            O => \N__29540\,
            I => \N__29529\
        );

    \I__7122\ : InMux
    port map (
            O => \N__29539\,
            I => \N__29526\
        );

    \I__7121\ : LocalMux
    port map (
            O => \N__29536\,
            I => \N__29521\
        );

    \I__7120\ : Span4Mux_h
    port map (
            O => \N__29533\,
            I => \N__29521\
        );

    \I__7119\ : InMux
    port map (
            O => \N__29532\,
            I => \N__29518\
        );

    \I__7118\ : LocalMux
    port map (
            O => \N__29529\,
            I => \N__29513\
        );

    \I__7117\ : LocalMux
    port map (
            O => \N__29526\,
            I => \N__29513\
        );

    \I__7116\ : Span4Mux_v
    port map (
            O => \N__29521\,
            I => \N__29509\
        );

    \I__7115\ : LocalMux
    port map (
            O => \N__29518\,
            I => \N__29506\
        );

    \I__7114\ : Span4Mux_v
    port map (
            O => \N__29513\,
            I => \N__29503\
        );

    \I__7113\ : InMux
    port map (
            O => \N__29512\,
            I => \N__29500\
        );

    \I__7112\ : Odrv4
    port map (
            O => \N__29509\,
            I => \Lab_UT.alarm_off\
        );

    \I__7111\ : Odrv12
    port map (
            O => \N__29506\,
            I => \Lab_UT.alarm_off\
        );

    \I__7110\ : Odrv4
    port map (
            O => \N__29503\,
            I => \Lab_UT.alarm_off\
        );

    \I__7109\ : LocalMux
    port map (
            O => \N__29500\,
            I => \Lab_UT.alarm_off\
        );

    \I__7108\ : CascadeMux
    port map (
            O => \N__29491\,
            I => \N__29487\
        );

    \I__7107\ : InMux
    port map (
            O => \N__29490\,
            I => \N__29484\
        );

    \I__7106\ : InMux
    port map (
            O => \N__29487\,
            I => \N__29481\
        );

    \I__7105\ : LocalMux
    port map (
            O => \N__29484\,
            I => \N__29367\
        );

    \I__7104\ : LocalMux
    port map (
            O => \N__29481\,
            I => \N__29364\
        );

    \I__7103\ : ClkMux
    port map (
            O => \N__29480\,
            I => \N__29137\
        );

    \I__7102\ : ClkMux
    port map (
            O => \N__29479\,
            I => \N__29137\
        );

    \I__7101\ : ClkMux
    port map (
            O => \N__29478\,
            I => \N__29137\
        );

    \I__7100\ : ClkMux
    port map (
            O => \N__29477\,
            I => \N__29137\
        );

    \I__7099\ : ClkMux
    port map (
            O => \N__29476\,
            I => \N__29137\
        );

    \I__7098\ : ClkMux
    port map (
            O => \N__29475\,
            I => \N__29137\
        );

    \I__7097\ : ClkMux
    port map (
            O => \N__29474\,
            I => \N__29137\
        );

    \I__7096\ : ClkMux
    port map (
            O => \N__29473\,
            I => \N__29137\
        );

    \I__7095\ : ClkMux
    port map (
            O => \N__29472\,
            I => \N__29137\
        );

    \I__7094\ : ClkMux
    port map (
            O => \N__29471\,
            I => \N__29137\
        );

    \I__7093\ : ClkMux
    port map (
            O => \N__29470\,
            I => \N__29137\
        );

    \I__7092\ : ClkMux
    port map (
            O => \N__29469\,
            I => \N__29137\
        );

    \I__7091\ : ClkMux
    port map (
            O => \N__29468\,
            I => \N__29137\
        );

    \I__7090\ : ClkMux
    port map (
            O => \N__29467\,
            I => \N__29137\
        );

    \I__7089\ : ClkMux
    port map (
            O => \N__29466\,
            I => \N__29137\
        );

    \I__7088\ : ClkMux
    port map (
            O => \N__29465\,
            I => \N__29137\
        );

    \I__7087\ : ClkMux
    port map (
            O => \N__29464\,
            I => \N__29137\
        );

    \I__7086\ : ClkMux
    port map (
            O => \N__29463\,
            I => \N__29137\
        );

    \I__7085\ : ClkMux
    port map (
            O => \N__29462\,
            I => \N__29137\
        );

    \I__7084\ : ClkMux
    port map (
            O => \N__29461\,
            I => \N__29137\
        );

    \I__7083\ : ClkMux
    port map (
            O => \N__29460\,
            I => \N__29137\
        );

    \I__7082\ : ClkMux
    port map (
            O => \N__29459\,
            I => \N__29137\
        );

    \I__7081\ : ClkMux
    port map (
            O => \N__29458\,
            I => \N__29137\
        );

    \I__7080\ : ClkMux
    port map (
            O => \N__29457\,
            I => \N__29137\
        );

    \I__7079\ : ClkMux
    port map (
            O => \N__29456\,
            I => \N__29137\
        );

    \I__7078\ : ClkMux
    port map (
            O => \N__29455\,
            I => \N__29137\
        );

    \I__7077\ : ClkMux
    port map (
            O => \N__29454\,
            I => \N__29137\
        );

    \I__7076\ : ClkMux
    port map (
            O => \N__29453\,
            I => \N__29137\
        );

    \I__7075\ : ClkMux
    port map (
            O => \N__29452\,
            I => \N__29137\
        );

    \I__7074\ : ClkMux
    port map (
            O => \N__29451\,
            I => \N__29137\
        );

    \I__7073\ : ClkMux
    port map (
            O => \N__29450\,
            I => \N__29137\
        );

    \I__7072\ : ClkMux
    port map (
            O => \N__29449\,
            I => \N__29137\
        );

    \I__7071\ : ClkMux
    port map (
            O => \N__29448\,
            I => \N__29137\
        );

    \I__7070\ : ClkMux
    port map (
            O => \N__29447\,
            I => \N__29137\
        );

    \I__7069\ : ClkMux
    port map (
            O => \N__29446\,
            I => \N__29137\
        );

    \I__7068\ : ClkMux
    port map (
            O => \N__29445\,
            I => \N__29137\
        );

    \I__7067\ : ClkMux
    port map (
            O => \N__29444\,
            I => \N__29137\
        );

    \I__7066\ : ClkMux
    port map (
            O => \N__29443\,
            I => \N__29137\
        );

    \I__7065\ : ClkMux
    port map (
            O => \N__29442\,
            I => \N__29137\
        );

    \I__7064\ : ClkMux
    port map (
            O => \N__29441\,
            I => \N__29137\
        );

    \I__7063\ : ClkMux
    port map (
            O => \N__29440\,
            I => \N__29137\
        );

    \I__7062\ : ClkMux
    port map (
            O => \N__29439\,
            I => \N__29137\
        );

    \I__7061\ : ClkMux
    port map (
            O => \N__29438\,
            I => \N__29137\
        );

    \I__7060\ : ClkMux
    port map (
            O => \N__29437\,
            I => \N__29137\
        );

    \I__7059\ : ClkMux
    port map (
            O => \N__29436\,
            I => \N__29137\
        );

    \I__7058\ : ClkMux
    port map (
            O => \N__29435\,
            I => \N__29137\
        );

    \I__7057\ : ClkMux
    port map (
            O => \N__29434\,
            I => \N__29137\
        );

    \I__7056\ : ClkMux
    port map (
            O => \N__29433\,
            I => \N__29137\
        );

    \I__7055\ : ClkMux
    port map (
            O => \N__29432\,
            I => \N__29137\
        );

    \I__7054\ : ClkMux
    port map (
            O => \N__29431\,
            I => \N__29137\
        );

    \I__7053\ : ClkMux
    port map (
            O => \N__29430\,
            I => \N__29137\
        );

    \I__7052\ : ClkMux
    port map (
            O => \N__29429\,
            I => \N__29137\
        );

    \I__7051\ : ClkMux
    port map (
            O => \N__29428\,
            I => \N__29137\
        );

    \I__7050\ : ClkMux
    port map (
            O => \N__29427\,
            I => \N__29137\
        );

    \I__7049\ : ClkMux
    port map (
            O => \N__29426\,
            I => \N__29137\
        );

    \I__7048\ : ClkMux
    port map (
            O => \N__29425\,
            I => \N__29137\
        );

    \I__7047\ : ClkMux
    port map (
            O => \N__29424\,
            I => \N__29137\
        );

    \I__7046\ : ClkMux
    port map (
            O => \N__29423\,
            I => \N__29137\
        );

    \I__7045\ : ClkMux
    port map (
            O => \N__29422\,
            I => \N__29137\
        );

    \I__7044\ : ClkMux
    port map (
            O => \N__29421\,
            I => \N__29137\
        );

    \I__7043\ : ClkMux
    port map (
            O => \N__29420\,
            I => \N__29137\
        );

    \I__7042\ : ClkMux
    port map (
            O => \N__29419\,
            I => \N__29137\
        );

    \I__7041\ : ClkMux
    port map (
            O => \N__29418\,
            I => \N__29137\
        );

    \I__7040\ : ClkMux
    port map (
            O => \N__29417\,
            I => \N__29137\
        );

    \I__7039\ : ClkMux
    port map (
            O => \N__29416\,
            I => \N__29137\
        );

    \I__7038\ : ClkMux
    port map (
            O => \N__29415\,
            I => \N__29137\
        );

    \I__7037\ : ClkMux
    port map (
            O => \N__29414\,
            I => \N__29137\
        );

    \I__7036\ : ClkMux
    port map (
            O => \N__29413\,
            I => \N__29137\
        );

    \I__7035\ : ClkMux
    port map (
            O => \N__29412\,
            I => \N__29137\
        );

    \I__7034\ : ClkMux
    port map (
            O => \N__29411\,
            I => \N__29137\
        );

    \I__7033\ : ClkMux
    port map (
            O => \N__29410\,
            I => \N__29137\
        );

    \I__7032\ : ClkMux
    port map (
            O => \N__29409\,
            I => \N__29137\
        );

    \I__7031\ : ClkMux
    port map (
            O => \N__29408\,
            I => \N__29137\
        );

    \I__7030\ : ClkMux
    port map (
            O => \N__29407\,
            I => \N__29137\
        );

    \I__7029\ : ClkMux
    port map (
            O => \N__29406\,
            I => \N__29137\
        );

    \I__7028\ : ClkMux
    port map (
            O => \N__29405\,
            I => \N__29137\
        );

    \I__7027\ : ClkMux
    port map (
            O => \N__29404\,
            I => \N__29137\
        );

    \I__7026\ : ClkMux
    port map (
            O => \N__29403\,
            I => \N__29137\
        );

    \I__7025\ : ClkMux
    port map (
            O => \N__29402\,
            I => \N__29137\
        );

    \I__7024\ : ClkMux
    port map (
            O => \N__29401\,
            I => \N__29137\
        );

    \I__7023\ : ClkMux
    port map (
            O => \N__29400\,
            I => \N__29137\
        );

    \I__7022\ : ClkMux
    port map (
            O => \N__29399\,
            I => \N__29137\
        );

    \I__7021\ : ClkMux
    port map (
            O => \N__29398\,
            I => \N__29137\
        );

    \I__7020\ : ClkMux
    port map (
            O => \N__29397\,
            I => \N__29137\
        );

    \I__7019\ : ClkMux
    port map (
            O => \N__29396\,
            I => \N__29137\
        );

    \I__7018\ : ClkMux
    port map (
            O => \N__29395\,
            I => \N__29137\
        );

    \I__7017\ : ClkMux
    port map (
            O => \N__29394\,
            I => \N__29137\
        );

    \I__7016\ : ClkMux
    port map (
            O => \N__29393\,
            I => \N__29137\
        );

    \I__7015\ : ClkMux
    port map (
            O => \N__29392\,
            I => \N__29137\
        );

    \I__7014\ : ClkMux
    port map (
            O => \N__29391\,
            I => \N__29137\
        );

    \I__7013\ : ClkMux
    port map (
            O => \N__29390\,
            I => \N__29137\
        );

    \I__7012\ : ClkMux
    port map (
            O => \N__29389\,
            I => \N__29137\
        );

    \I__7011\ : ClkMux
    port map (
            O => \N__29388\,
            I => \N__29137\
        );

    \I__7010\ : ClkMux
    port map (
            O => \N__29387\,
            I => \N__29137\
        );

    \I__7009\ : ClkMux
    port map (
            O => \N__29386\,
            I => \N__29137\
        );

    \I__7008\ : ClkMux
    port map (
            O => \N__29385\,
            I => \N__29137\
        );

    \I__7007\ : ClkMux
    port map (
            O => \N__29384\,
            I => \N__29137\
        );

    \I__7006\ : ClkMux
    port map (
            O => \N__29383\,
            I => \N__29137\
        );

    \I__7005\ : ClkMux
    port map (
            O => \N__29382\,
            I => \N__29137\
        );

    \I__7004\ : ClkMux
    port map (
            O => \N__29381\,
            I => \N__29137\
        );

    \I__7003\ : ClkMux
    port map (
            O => \N__29380\,
            I => \N__29137\
        );

    \I__7002\ : ClkMux
    port map (
            O => \N__29379\,
            I => \N__29137\
        );

    \I__7001\ : ClkMux
    port map (
            O => \N__29378\,
            I => \N__29137\
        );

    \I__7000\ : ClkMux
    port map (
            O => \N__29377\,
            I => \N__29137\
        );

    \I__6999\ : ClkMux
    port map (
            O => \N__29376\,
            I => \N__29137\
        );

    \I__6998\ : ClkMux
    port map (
            O => \N__29375\,
            I => \N__29137\
        );

    \I__6997\ : ClkMux
    port map (
            O => \N__29374\,
            I => \N__29137\
        );

    \I__6996\ : ClkMux
    port map (
            O => \N__29373\,
            I => \N__29137\
        );

    \I__6995\ : ClkMux
    port map (
            O => \N__29372\,
            I => \N__29137\
        );

    \I__6994\ : ClkMux
    port map (
            O => \N__29371\,
            I => \N__29137\
        );

    \I__6993\ : ClkMux
    port map (
            O => \N__29370\,
            I => \N__29137\
        );

    \I__6992\ : Glb2LocalMux
    port map (
            O => \N__29367\,
            I => \N__29137\
        );

    \I__6991\ : Glb2LocalMux
    port map (
            O => \N__29364\,
            I => \N__29137\
        );

    \I__6990\ : GlobalMux
    port map (
            O => \N__29137\,
            I => \N__29134\
        );

    \I__6989\ : gio2CtrlBuf
    port map (
            O => \N__29134\,
            I => clk_g
        );

    \I__6988\ : SRMux
    port map (
            O => \N__29131\,
            I => \N__29127\
        );

    \I__6987\ : CascadeMux
    port map (
            O => \N__29130\,
            I => \N__29123\
        );

    \I__6986\ : LocalMux
    port map (
            O => \N__29127\,
            I => \N__29120\
        );

    \I__6985\ : InMux
    port map (
            O => \N__29126\,
            I => \N__29115\
        );

    \I__6984\ : InMux
    port map (
            O => \N__29123\,
            I => \N__29115\
        );

    \I__6983\ : Odrv12
    port map (
            O => \N__29120\,
            I => \Lab_UT.dictrl.nextState_al22\
        );

    \I__6982\ : LocalMux
    port map (
            O => \N__29115\,
            I => \Lab_UT.dictrl.nextState_al22\
        );

    \I__6981\ : CascadeMux
    port map (
            O => \N__29110\,
            I => \Lab_UT.didp.Mones_subtractor.un1_q_axb_0_cascade_\
        );

    \I__6980\ : InMux
    port map (
            O => \N__29107\,
            I => \N__29099\
        );

    \I__6979\ : CascadeMux
    port map (
            O => \N__29106\,
            I => \N__29094\
        );

    \I__6978\ : InMux
    port map (
            O => \N__29105\,
            I => \N__29091\
        );

    \I__6977\ : InMux
    port map (
            O => \N__29104\,
            I => \N__29086\
        );

    \I__6976\ : InMux
    port map (
            O => \N__29103\,
            I => \N__29086\
        );

    \I__6975\ : InMux
    port map (
            O => \N__29102\,
            I => \N__29083\
        );

    \I__6974\ : LocalMux
    port map (
            O => \N__29099\,
            I => \N__29080\
        );

    \I__6973\ : InMux
    port map (
            O => \N__29098\,
            I => \N__29077\
        );

    \I__6972\ : InMux
    port map (
            O => \N__29097\,
            I => \N__29074\
        );

    \I__6971\ : InMux
    port map (
            O => \N__29094\,
            I => \N__29070\
        );

    \I__6970\ : LocalMux
    port map (
            O => \N__29091\,
            I => \N__29065\
        );

    \I__6969\ : LocalMux
    port map (
            O => \N__29086\,
            I => \N__29065\
        );

    \I__6968\ : LocalMux
    port map (
            O => \N__29083\,
            I => \N__29059\
        );

    \I__6967\ : Span4Mux_s0_h
    port map (
            O => \N__29080\,
            I => \N__29052\
        );

    \I__6966\ : LocalMux
    port map (
            O => \N__29077\,
            I => \N__29052\
        );

    \I__6965\ : LocalMux
    port map (
            O => \N__29074\,
            I => \N__29052\
        );

    \I__6964\ : InMux
    port map (
            O => \N__29073\,
            I => \N__29049\
        );

    \I__6963\ : LocalMux
    port map (
            O => \N__29070\,
            I => \N__29042\
        );

    \I__6962\ : Span4Mux_v
    port map (
            O => \N__29065\,
            I => \N__29042\
        );

    \I__6961\ : InMux
    port map (
            O => \N__29064\,
            I => \N__29035\
        );

    \I__6960\ : InMux
    port map (
            O => \N__29063\,
            I => \N__29035\
        );

    \I__6959\ : InMux
    port map (
            O => \N__29062\,
            I => \N__29035\
        );

    \I__6958\ : Span4Mux_v
    port map (
            O => \N__29059\,
            I => \N__29030\
        );

    \I__6957\ : Span4Mux_v
    port map (
            O => \N__29052\,
            I => \N__29030\
        );

    \I__6956\ : LocalMux
    port map (
            O => \N__29049\,
            I => \N__29027\
        );

    \I__6955\ : CascadeMux
    port map (
            O => \N__29048\,
            I => \N__29023\
        );

    \I__6954\ : CascadeMux
    port map (
            O => \N__29047\,
            I => \N__29020\
        );

    \I__6953\ : Span4Mux_v
    port map (
            O => \N__29042\,
            I => \N__29015\
        );

    \I__6952\ : LocalMux
    port map (
            O => \N__29035\,
            I => \N__29015\
        );

    \I__6951\ : Span4Mux_h
    port map (
            O => \N__29030\,
            I => \N__29010\
        );

    \I__6950\ : Span4Mux_h
    port map (
            O => \N__29027\,
            I => \N__29010\
        );

    \I__6949\ : InMux
    port map (
            O => \N__29026\,
            I => \N__29003\
        );

    \I__6948\ : InMux
    port map (
            O => \N__29023\,
            I => \N__29003\
        );

    \I__6947\ : InMux
    port map (
            O => \N__29020\,
            I => \N__29003\
        );

    \I__6946\ : Odrv4
    port map (
            O => \N__29015\,
            I => bu_rx_data_0
        );

    \I__6945\ : Odrv4
    port map (
            O => \N__29010\,
            I => bu_rx_data_0
        );

    \I__6944\ : LocalMux
    port map (
            O => \N__29003\,
            I => bu_rx_data_0
        );

    \I__6943\ : InMux
    port map (
            O => \N__28996\,
            I => \N__28991\
        );

    \I__6942\ : CascadeMux
    port map (
            O => \N__28995\,
            I => \N__28988\
        );

    \I__6941\ : CascadeMux
    port map (
            O => \N__28994\,
            I => \N__28975\
        );

    \I__6940\ : LocalMux
    port map (
            O => \N__28991\,
            I => \N__28971\
        );

    \I__6939\ : InMux
    port map (
            O => \N__28988\,
            I => \N__28968\
        );

    \I__6938\ : InMux
    port map (
            O => \N__28987\,
            I => \N__28965\
        );

    \I__6937\ : InMux
    port map (
            O => \N__28986\,
            I => \N__28957\
        );

    \I__6936\ : InMux
    port map (
            O => \N__28985\,
            I => \N__28957\
        );

    \I__6935\ : InMux
    port map (
            O => \N__28984\,
            I => \N__28957\
        );

    \I__6934\ : InMux
    port map (
            O => \N__28983\,
            I => \N__28954\
        );

    \I__6933\ : InMux
    port map (
            O => \N__28982\,
            I => \N__28951\
        );

    \I__6932\ : InMux
    port map (
            O => \N__28981\,
            I => \N__28948\
        );

    \I__6931\ : InMux
    port map (
            O => \N__28980\,
            I => \N__28944\
        );

    \I__6930\ : InMux
    port map (
            O => \N__28979\,
            I => \N__28938\
        );

    \I__6929\ : InMux
    port map (
            O => \N__28978\,
            I => \N__28938\
        );

    \I__6928\ : InMux
    port map (
            O => \N__28975\,
            I => \N__28935\
        );

    \I__6927\ : InMux
    port map (
            O => \N__28974\,
            I => \N__28932\
        );

    \I__6926\ : Span4Mux_v
    port map (
            O => \N__28971\,
            I => \N__28925\
        );

    \I__6925\ : LocalMux
    port map (
            O => \N__28968\,
            I => \N__28925\
        );

    \I__6924\ : LocalMux
    port map (
            O => \N__28965\,
            I => \N__28925\
        );

    \I__6923\ : CascadeMux
    port map (
            O => \N__28964\,
            I => \N__28921\
        );

    \I__6922\ : LocalMux
    port map (
            O => \N__28957\,
            I => \N__28916\
        );

    \I__6921\ : LocalMux
    port map (
            O => \N__28954\,
            I => \N__28916\
        );

    \I__6920\ : LocalMux
    port map (
            O => \N__28951\,
            I => \N__28913\
        );

    \I__6919\ : LocalMux
    port map (
            O => \N__28948\,
            I => \N__28910\
        );

    \I__6918\ : CascadeMux
    port map (
            O => \N__28947\,
            I => \N__28907\
        );

    \I__6917\ : LocalMux
    port map (
            O => \N__28944\,
            I => \N__28902\
        );

    \I__6916\ : CascadeMux
    port map (
            O => \N__28943\,
            I => \N__28899\
        );

    \I__6915\ : LocalMux
    port map (
            O => \N__28938\,
            I => \N__28896\
        );

    \I__6914\ : LocalMux
    port map (
            O => \N__28935\,
            I => \N__28893\
        );

    \I__6913\ : LocalMux
    port map (
            O => \N__28932\,
            I => \N__28890\
        );

    \I__6912\ : Span4Mux_h
    port map (
            O => \N__28925\,
            I => \N__28887\
        );

    \I__6911\ : InMux
    port map (
            O => \N__28924\,
            I => \N__28884\
        );

    \I__6910\ : InMux
    port map (
            O => \N__28921\,
            I => \N__28881\
        );

    \I__6909\ : Span4Mux_v
    port map (
            O => \N__28916\,
            I => \N__28878\
        );

    \I__6908\ : Span4Mux_v
    port map (
            O => \N__28913\,
            I => \N__28873\
        );

    \I__6907\ : Span4Mux_h
    port map (
            O => \N__28910\,
            I => \N__28873\
        );

    \I__6906\ : InMux
    port map (
            O => \N__28907\,
            I => \N__28870\
        );

    \I__6905\ : InMux
    port map (
            O => \N__28906\,
            I => \N__28867\
        );

    \I__6904\ : InMux
    port map (
            O => \N__28905\,
            I => \N__28864\
        );

    \I__6903\ : Span12Mux_v
    port map (
            O => \N__28902\,
            I => \N__28861\
        );

    \I__6902\ : InMux
    port map (
            O => \N__28899\,
            I => \N__28858\
        );

    \I__6901\ : Span4Mux_v
    port map (
            O => \N__28896\,
            I => \N__28851\
        );

    \I__6900\ : Span4Mux_v
    port map (
            O => \N__28893\,
            I => \N__28851\
        );

    \I__6899\ : Span4Mux_s1_v
    port map (
            O => \N__28890\,
            I => \N__28851\
        );

    \I__6898\ : Span4Mux_v
    port map (
            O => \N__28887\,
            I => \N__28844\
        );

    \I__6897\ : LocalMux
    port map (
            O => \N__28884\,
            I => \N__28844\
        );

    \I__6896\ : LocalMux
    port map (
            O => \N__28881\,
            I => \N__28844\
        );

    \I__6895\ : Span4Mux_v
    port map (
            O => \N__28878\,
            I => \N__28837\
        );

    \I__6894\ : Span4Mux_h
    port map (
            O => \N__28873\,
            I => \N__28837\
        );

    \I__6893\ : LocalMux
    port map (
            O => \N__28870\,
            I => \N__28837\
        );

    \I__6892\ : LocalMux
    port map (
            O => \N__28867\,
            I => bu_rx_data_3
        );

    \I__6891\ : LocalMux
    port map (
            O => \N__28864\,
            I => bu_rx_data_3
        );

    \I__6890\ : Odrv12
    port map (
            O => \N__28861\,
            I => bu_rx_data_3
        );

    \I__6889\ : LocalMux
    port map (
            O => \N__28858\,
            I => bu_rx_data_3
        );

    \I__6888\ : Odrv4
    port map (
            O => \N__28851\,
            I => bu_rx_data_3
        );

    \I__6887\ : Odrv4
    port map (
            O => \N__28844\,
            I => bu_rx_data_3
        );

    \I__6886\ : Odrv4
    port map (
            O => \N__28837\,
            I => bu_rx_data_3
        );

    \I__6885\ : CascadeMux
    port map (
            O => \N__28822\,
            I => \N__28813\
        );

    \I__6884\ : InMux
    port map (
            O => \N__28821\,
            I => \N__28809\
        );

    \I__6883\ : InMux
    port map (
            O => \N__28820\,
            I => \N__28806\
        );

    \I__6882\ : InMux
    port map (
            O => \N__28819\,
            I => \N__28803\
        );

    \I__6881\ : InMux
    port map (
            O => \N__28818\,
            I => \N__28800\
        );

    \I__6880\ : InMux
    port map (
            O => \N__28817\,
            I => \N__28797\
        );

    \I__6879\ : InMux
    port map (
            O => \N__28816\,
            I => \N__28792\
        );

    \I__6878\ : InMux
    port map (
            O => \N__28813\,
            I => \N__28789\
        );

    \I__6877\ : InMux
    port map (
            O => \N__28812\,
            I => \N__28786\
        );

    \I__6876\ : LocalMux
    port map (
            O => \N__28809\,
            I => \N__28783\
        );

    \I__6875\ : LocalMux
    port map (
            O => \N__28806\,
            I => \N__28776\
        );

    \I__6874\ : LocalMux
    port map (
            O => \N__28803\,
            I => \N__28776\
        );

    \I__6873\ : LocalMux
    port map (
            O => \N__28800\,
            I => \N__28776\
        );

    \I__6872\ : LocalMux
    port map (
            O => \N__28797\,
            I => \N__28773\
        );

    \I__6871\ : InMux
    port map (
            O => \N__28796\,
            I => \N__28766\
        );

    \I__6870\ : InMux
    port map (
            O => \N__28795\,
            I => \N__28766\
        );

    \I__6869\ : LocalMux
    port map (
            O => \N__28792\,
            I => \N__28763\
        );

    \I__6868\ : LocalMux
    port map (
            O => \N__28789\,
            I => \N__28760\
        );

    \I__6867\ : LocalMux
    port map (
            O => \N__28786\,
            I => \N__28757\
        );

    \I__6866\ : Span4Mux_v
    port map (
            O => \N__28783\,
            I => \N__28750\
        );

    \I__6865\ : Span4Mux_v
    port map (
            O => \N__28776\,
            I => \N__28747\
        );

    \I__6864\ : Span4Mux_s2_v
    port map (
            O => \N__28773\,
            I => \N__28744\
        );

    \I__6863\ : InMux
    port map (
            O => \N__28772\,
            I => \N__28738\
        );

    \I__6862\ : InMux
    port map (
            O => \N__28771\,
            I => \N__28738\
        );

    \I__6861\ : LocalMux
    port map (
            O => \N__28766\,
            I => \N__28735\
        );

    \I__6860\ : Span4Mux_v
    port map (
            O => \N__28763\,
            I => \N__28732\
        );

    \I__6859\ : Span4Mux_s2_h
    port map (
            O => \N__28760\,
            I => \N__28729\
        );

    \I__6858\ : Span12Mux_s8_h
    port map (
            O => \N__28757\,
            I => \N__28726\
        );

    \I__6857\ : InMux
    port map (
            O => \N__28756\,
            I => \N__28721\
        );

    \I__6856\ : InMux
    port map (
            O => \N__28755\,
            I => \N__28721\
        );

    \I__6855\ : InMux
    port map (
            O => \N__28754\,
            I => \N__28718\
        );

    \I__6854\ : InMux
    port map (
            O => \N__28753\,
            I => \N__28715\
        );

    \I__6853\ : Span4Mux_v
    port map (
            O => \N__28750\,
            I => \N__28708\
        );

    \I__6852\ : Span4Mux_v
    port map (
            O => \N__28747\,
            I => \N__28708\
        );

    \I__6851\ : Span4Mux_h
    port map (
            O => \N__28744\,
            I => \N__28708\
        );

    \I__6850\ : InMux
    port map (
            O => \N__28743\,
            I => \N__28705\
        );

    \I__6849\ : LocalMux
    port map (
            O => \N__28738\,
            I => bu_rx_data_1
        );

    \I__6848\ : Odrv12
    port map (
            O => \N__28735\,
            I => bu_rx_data_1
        );

    \I__6847\ : Odrv4
    port map (
            O => \N__28732\,
            I => bu_rx_data_1
        );

    \I__6846\ : Odrv4
    port map (
            O => \N__28729\,
            I => bu_rx_data_1
        );

    \I__6845\ : Odrv12
    port map (
            O => \N__28726\,
            I => bu_rx_data_1
        );

    \I__6844\ : LocalMux
    port map (
            O => \N__28721\,
            I => bu_rx_data_1
        );

    \I__6843\ : LocalMux
    port map (
            O => \N__28718\,
            I => bu_rx_data_1
        );

    \I__6842\ : LocalMux
    port map (
            O => \N__28715\,
            I => bu_rx_data_1
        );

    \I__6841\ : Odrv4
    port map (
            O => \N__28708\,
            I => bu_rx_data_1
        );

    \I__6840\ : LocalMux
    port map (
            O => \N__28705\,
            I => bu_rx_data_1
        );

    \I__6839\ : InMux
    port map (
            O => \N__28684\,
            I => \N__28679\
        );

    \I__6838\ : InMux
    port map (
            O => \N__28683\,
            I => \N__28672\
        );

    \I__6837\ : InMux
    port map (
            O => \N__28682\,
            I => \N__28672\
        );

    \I__6836\ : LocalMux
    port map (
            O => \N__28679\,
            I => \N__28669\
        );

    \I__6835\ : InMux
    port map (
            O => \N__28678\,
            I => \N__28666\
        );

    \I__6834\ : CascadeMux
    port map (
            O => \N__28677\,
            I => \N__28661\
        );

    \I__6833\ : LocalMux
    port map (
            O => \N__28672\,
            I => \N__28653\
        );

    \I__6832\ : Span4Mux_v
    port map (
            O => \N__28669\,
            I => \N__28653\
        );

    \I__6831\ : LocalMux
    port map (
            O => \N__28666\,
            I => \N__28653\
        );

    \I__6830\ : InMux
    port map (
            O => \N__28665\,
            I => \N__28644\
        );

    \I__6829\ : InMux
    port map (
            O => \N__28664\,
            I => \N__28644\
        );

    \I__6828\ : InMux
    port map (
            O => \N__28661\,
            I => \N__28644\
        );

    \I__6827\ : InMux
    port map (
            O => \N__28660\,
            I => \N__28644\
        );

    \I__6826\ : Span4Mux_v
    port map (
            O => \N__28653\,
            I => \N__28641\
        );

    \I__6825\ : LocalMux
    port map (
            O => \N__28644\,
            I => \Lab_UT.didp.N_84\
        );

    \I__6824\ : Odrv4
    port map (
            O => \N__28641\,
            I => \Lab_UT.didp.N_84\
        );

    \I__6823\ : InMux
    port map (
            O => \N__28636\,
            I => \N__28624\
        );

    \I__6822\ : InMux
    port map (
            O => \N__28635\,
            I => \N__28624\
        );

    \I__6821\ : InMux
    port map (
            O => \N__28634\,
            I => \N__28624\
        );

    \I__6820\ : InMux
    port map (
            O => \N__28633\,
            I => \N__28624\
        );

    \I__6819\ : LocalMux
    port map (
            O => \N__28624\,
            I => \N__28621\
        );

    \I__6818\ : Odrv4
    port map (
            O => \N__28621\,
            I => \Lab_UT.didp.Mones_subtractor.q_0_sqmuxa\
        );

    \I__6817\ : CascadeMux
    port map (
            O => \N__28618\,
            I => \Lab_UT.didp.Mones_subtractor.q_RNO_0_2_2_cascade_\
        );

    \I__6816\ : InMux
    port map (
            O => \N__28615\,
            I => \N__28603\
        );

    \I__6815\ : InMux
    port map (
            O => \N__28614\,
            I => \N__28598\
        );

    \I__6814\ : InMux
    port map (
            O => \N__28613\,
            I => \N__28593\
        );

    \I__6813\ : CascadeMux
    port map (
            O => \N__28612\,
            I => \N__28590\
        );

    \I__6812\ : InMux
    port map (
            O => \N__28611\,
            I => \N__28585\
        );

    \I__6811\ : InMux
    port map (
            O => \N__28610\,
            I => \N__28585\
        );

    \I__6810\ : InMux
    port map (
            O => \N__28609\,
            I => \N__28580\
        );

    \I__6809\ : InMux
    port map (
            O => \N__28608\,
            I => \N__28580\
        );

    \I__6808\ : InMux
    port map (
            O => \N__28607\,
            I => \N__28577\
        );

    \I__6807\ : InMux
    port map (
            O => \N__28606\,
            I => \N__28574\
        );

    \I__6806\ : LocalMux
    port map (
            O => \N__28603\,
            I => \N__28570\
        );

    \I__6805\ : InMux
    port map (
            O => \N__28602\,
            I => \N__28567\
        );

    \I__6804\ : InMux
    port map (
            O => \N__28601\,
            I => \N__28564\
        );

    \I__6803\ : LocalMux
    port map (
            O => \N__28598\,
            I => \N__28560\
        );

    \I__6802\ : InMux
    port map (
            O => \N__28597\,
            I => \N__28557\
        );

    \I__6801\ : InMux
    port map (
            O => \N__28596\,
            I => \N__28554\
        );

    \I__6800\ : LocalMux
    port map (
            O => \N__28593\,
            I => \N__28551\
        );

    \I__6799\ : InMux
    port map (
            O => \N__28590\,
            I => \N__28548\
        );

    \I__6798\ : LocalMux
    port map (
            O => \N__28585\,
            I => \N__28543\
        );

    \I__6797\ : LocalMux
    port map (
            O => \N__28580\,
            I => \N__28543\
        );

    \I__6796\ : LocalMux
    port map (
            O => \N__28577\,
            I => \N__28540\
        );

    \I__6795\ : LocalMux
    port map (
            O => \N__28574\,
            I => \N__28536\
        );

    \I__6794\ : InMux
    port map (
            O => \N__28573\,
            I => \N__28533\
        );

    \I__6793\ : Span4Mux_v
    port map (
            O => \N__28570\,
            I => \N__28530\
        );

    \I__6792\ : LocalMux
    port map (
            O => \N__28567\,
            I => \N__28527\
        );

    \I__6791\ : LocalMux
    port map (
            O => \N__28564\,
            I => \N__28524\
        );

    \I__6790\ : InMux
    port map (
            O => \N__28563\,
            I => \N__28521\
        );

    \I__6789\ : Span4Mux_v
    port map (
            O => \N__28560\,
            I => \N__28518\
        );

    \I__6788\ : LocalMux
    port map (
            O => \N__28557\,
            I => \N__28515\
        );

    \I__6787\ : LocalMux
    port map (
            O => \N__28554\,
            I => \N__28510\
        );

    \I__6786\ : Span4Mux_s2_v
    port map (
            O => \N__28551\,
            I => \N__28510\
        );

    \I__6785\ : LocalMux
    port map (
            O => \N__28548\,
            I => \N__28500\
        );

    \I__6784\ : Span12Mux_s7_v
    port map (
            O => \N__28543\,
            I => \N__28500\
        );

    \I__6783\ : Span12Mux_s3_h
    port map (
            O => \N__28540\,
            I => \N__28500\
        );

    \I__6782\ : InMux
    port map (
            O => \N__28539\,
            I => \N__28497\
        );

    \I__6781\ : Span4Mux_h
    port map (
            O => \N__28536\,
            I => \N__28494\
        );

    \I__6780\ : LocalMux
    port map (
            O => \N__28533\,
            I => \N__28485\
        );

    \I__6779\ : Span4Mux_v
    port map (
            O => \N__28530\,
            I => \N__28485\
        );

    \I__6778\ : Span4Mux_v
    port map (
            O => \N__28527\,
            I => \N__28485\
        );

    \I__6777\ : Span4Mux_s2_v
    port map (
            O => \N__28524\,
            I => \N__28485\
        );

    \I__6776\ : LocalMux
    port map (
            O => \N__28521\,
            I => \N__28476\
        );

    \I__6775\ : Span4Mux_v
    port map (
            O => \N__28518\,
            I => \N__28476\
        );

    \I__6774\ : Span4Mux_s2_v
    port map (
            O => \N__28515\,
            I => \N__28476\
        );

    \I__6773\ : Span4Mux_h
    port map (
            O => \N__28510\,
            I => \N__28476\
        );

    \I__6772\ : InMux
    port map (
            O => \N__28509\,
            I => \N__28469\
        );

    \I__6771\ : InMux
    port map (
            O => \N__28508\,
            I => \N__28469\
        );

    \I__6770\ : InMux
    port map (
            O => \N__28507\,
            I => \N__28469\
        );

    \I__6769\ : Odrv12
    port map (
            O => \N__28500\,
            I => bu_rx_data_2
        );

    \I__6768\ : LocalMux
    port map (
            O => \N__28497\,
            I => bu_rx_data_2
        );

    \I__6767\ : Odrv4
    port map (
            O => \N__28494\,
            I => bu_rx_data_2
        );

    \I__6766\ : Odrv4
    port map (
            O => \N__28485\,
            I => bu_rx_data_2
        );

    \I__6765\ : Odrv4
    port map (
            O => \N__28476\,
            I => bu_rx_data_2
        );

    \I__6764\ : LocalMux
    port map (
            O => \N__28469\,
            I => bu_rx_data_2
        );

    \I__6763\ : SRMux
    port map (
            O => \N__28456\,
            I => \N__28452\
        );

    \I__6762\ : SRMux
    port map (
            O => \N__28455\,
            I => \N__28449\
        );

    \I__6761\ : LocalMux
    port map (
            O => \N__28452\,
            I => \N__28443\
        );

    \I__6760\ : LocalMux
    port map (
            O => \N__28449\,
            I => \N__28440\
        );

    \I__6759\ : SRMux
    port map (
            O => \N__28448\,
            I => \N__28437\
        );

    \I__6758\ : SRMux
    port map (
            O => \N__28447\,
            I => \N__28433\
        );

    \I__6757\ : SRMux
    port map (
            O => \N__28446\,
            I => \N__28430\
        );

    \I__6756\ : Span4Mux_s3_h
    port map (
            O => \N__28443\,
            I => \N__28423\
        );

    \I__6755\ : Span4Mux_s3_h
    port map (
            O => \N__28440\,
            I => \N__28423\
        );

    \I__6754\ : LocalMux
    port map (
            O => \N__28437\,
            I => \N__28423\
        );

    \I__6753\ : SRMux
    port map (
            O => \N__28436\,
            I => \N__28420\
        );

    \I__6752\ : LocalMux
    port map (
            O => \N__28433\,
            I => \N__28416\
        );

    \I__6751\ : LocalMux
    port map (
            O => \N__28430\,
            I => \N__28413\
        );

    \I__6750\ : Span4Mux_v
    port map (
            O => \N__28423\,
            I => \N__28408\
        );

    \I__6749\ : LocalMux
    port map (
            O => \N__28420\,
            I => \N__28408\
        );

    \I__6748\ : SRMux
    port map (
            O => \N__28419\,
            I => \N__28405\
        );

    \I__6747\ : Span4Mux_v
    port map (
            O => \N__28416\,
            I => \N__28402\
        );

    \I__6746\ : Span4Mux_s3_h
    port map (
            O => \N__28413\,
            I => \N__28399\
        );

    \I__6745\ : Span4Mux_s3_h
    port map (
            O => \N__28408\,
            I => \N__28396\
        );

    \I__6744\ : LocalMux
    port map (
            O => \N__28405\,
            I => \N__28393\
        );

    \I__6743\ : Span4Mux_h
    port map (
            O => \N__28402\,
            I => \N__28390\
        );

    \I__6742\ : Span4Mux_h
    port map (
            O => \N__28399\,
            I => \N__28387\
        );

    \I__6741\ : Span4Mux_h
    port map (
            O => \N__28396\,
            I => \N__28384\
        );

    \I__6740\ : Span4Mux_s3_h
    port map (
            O => \N__28393\,
            I => \N__28381\
        );

    \I__6739\ : Span4Mux_h
    port map (
            O => \N__28390\,
            I => \N__28378\
        );

    \I__6738\ : Span4Mux_v
    port map (
            O => \N__28387\,
            I => \N__28375\
        );

    \I__6737\ : Span4Mux_v
    port map (
            O => \N__28384\,
            I => \N__28372\
        );

    \I__6736\ : Span4Mux_h
    port map (
            O => \N__28381\,
            I => \N__28369\
        );

    \I__6735\ : Odrv4
    port map (
            O => \N__28378\,
            I => \Lab_UT.didp.q20_0_i\
        );

    \I__6734\ : Odrv4
    port map (
            O => \N__28375\,
            I => \Lab_UT.didp.q20_0_i\
        );

    \I__6733\ : Odrv4
    port map (
            O => \N__28372\,
            I => \Lab_UT.didp.q20_0_i\
        );

    \I__6732\ : Odrv4
    port map (
            O => \N__28369\,
            I => \Lab_UT.didp.q20_0_i\
        );

    \I__6731\ : InMux
    port map (
            O => \N__28360\,
            I => \Lab_UT.didp.Mones_subtractor.un1_q_cry_0_s1\
        );

    \I__6730\ : CascadeMux
    port map (
            O => \N__28357\,
            I => \N__28350\
        );

    \I__6729\ : CascadeMux
    port map (
            O => \N__28356\,
            I => \N__28347\
        );

    \I__6728\ : SRMux
    port map (
            O => \N__28355\,
            I => \N__28344\
        );

    \I__6727\ : IoInMux
    port map (
            O => \N__28354\,
            I => \N__28341\
        );

    \I__6726\ : InMux
    port map (
            O => \N__28353\,
            I => \N__28336\
        );

    \I__6725\ : InMux
    port map (
            O => \N__28350\,
            I => \N__28336\
        );

    \I__6724\ : InMux
    port map (
            O => \N__28347\,
            I => \N__28333\
        );

    \I__6723\ : LocalMux
    port map (
            O => \N__28344\,
            I => \N__28330\
        );

    \I__6722\ : LocalMux
    port map (
            O => \N__28341\,
            I => \N__28327\
        );

    \I__6721\ : LocalMux
    port map (
            O => \N__28336\,
            I => \N__28324\
        );

    \I__6720\ : LocalMux
    port map (
            O => \N__28333\,
            I => \N__28321\
        );

    \I__6719\ : Span4Mux_h
    port map (
            O => \N__28330\,
            I => \N__28318\
        );

    \I__6718\ : Span4Mux_s3_v
    port map (
            O => \N__28327\,
            I => \N__28315\
        );

    \I__6717\ : Span12Mux_s6_h
    port map (
            O => \N__28324\,
            I => \N__28312\
        );

    \I__6716\ : Span12Mux_s11_v
    port map (
            O => \N__28321\,
            I => \N__28309\
        );

    \I__6715\ : Span4Mux_h
    port map (
            O => \N__28318\,
            I => \N__28304\
        );

    \I__6714\ : Span4Mux_h
    port map (
            O => \N__28315\,
            I => \N__28304\
        );

    \I__6713\ : Odrv12
    port map (
            O => \N__28312\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6712\ : Odrv12
    port map (
            O => \N__28309\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6711\ : Odrv4
    port map (
            O => \N__28304\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6710\ : InMux
    port map (
            O => \N__28297\,
            I => \N__28290\
        );

    \I__6709\ : InMux
    port map (
            O => \N__28296\,
            I => \N__28290\
        );

    \I__6708\ : CascadeMux
    port map (
            O => \N__28295\,
            I => \N__28287\
        );

    \I__6707\ : LocalMux
    port map (
            O => \N__28290\,
            I => \N__28282\
        );

    \I__6706\ : InMux
    port map (
            O => \N__28287\,
            I => \N__28279\
        );

    \I__6705\ : InMux
    port map (
            O => \N__28286\,
            I => \N__28274\
        );

    \I__6704\ : InMux
    port map (
            O => \N__28285\,
            I => \N__28274\
        );

    \I__6703\ : Sp12to4
    port map (
            O => \N__28282\,
            I => \N__28271\
        );

    \I__6702\ : LocalMux
    port map (
            O => \N__28279\,
            I => \Lab_UT.didp.di_Mones_2\
        );

    \I__6701\ : LocalMux
    port map (
            O => \N__28274\,
            I => \Lab_UT.didp.di_Mones_2\
        );

    \I__6700\ : Odrv12
    port map (
            O => \N__28271\,
            I => \Lab_UT.didp.di_Mones_2\
        );

    \I__6699\ : InMux
    port map (
            O => \N__28264\,
            I => \N__28261\
        );

    \I__6698\ : LocalMux
    port map (
            O => \N__28261\,
            I => \N__28258\
        );

    \I__6697\ : Odrv4
    port map (
            O => \N__28258\,
            I => \Lab_UT.didp.Mones_subtractor.un1_q_cry_1_s1_THRU_CO\
        );

    \I__6696\ : InMux
    port map (
            O => \N__28255\,
            I => \Lab_UT.didp.Mones_subtractor.un1_q_cry_1_s1\
        );

    \I__6695\ : InMux
    port map (
            O => \N__28252\,
            I => \N__28248\
        );

    \I__6694\ : InMux
    port map (
            O => \N__28251\,
            I => \N__28244\
        );

    \I__6693\ : LocalMux
    port map (
            O => \N__28248\,
            I => \N__28241\
        );

    \I__6692\ : CascadeMux
    port map (
            O => \N__28247\,
            I => \N__28237\
        );

    \I__6691\ : LocalMux
    port map (
            O => \N__28244\,
            I => \N__28234\
        );

    \I__6690\ : Span4Mux_h
    port map (
            O => \N__28241\,
            I => \N__28231\
        );

    \I__6689\ : InMux
    port map (
            O => \N__28240\,
            I => \N__28228\
        );

    \I__6688\ : InMux
    port map (
            O => \N__28237\,
            I => \N__28225\
        );

    \I__6687\ : Span4Mux_h
    port map (
            O => \N__28234\,
            I => \N__28222\
        );

    \I__6686\ : Odrv4
    port map (
            O => \N__28231\,
            I => \Lab_UT.didp.di_Mones_3\
        );

    \I__6685\ : LocalMux
    port map (
            O => \N__28228\,
            I => \Lab_UT.didp.di_Mones_3\
        );

    \I__6684\ : LocalMux
    port map (
            O => \N__28225\,
            I => \Lab_UT.didp.di_Mones_3\
        );

    \I__6683\ : Odrv4
    port map (
            O => \N__28222\,
            I => \Lab_UT.didp.di_Mones_3\
        );

    \I__6682\ : InMux
    port map (
            O => \N__28213\,
            I => \Lab_UT.didp.Mones_subtractor.un1_q_cry_2_s1\
        );

    \I__6681\ : CascadeMux
    port map (
            O => \N__28210\,
            I => \Lab_UT.ld_enable_Sones_cascade_\
        );

    \I__6680\ : InMux
    port map (
            O => \N__28207\,
            I => \N__28204\
        );

    \I__6679\ : LocalMux
    port map (
            O => \N__28204\,
            I => \Lab_UT.didp.Sones_subtractor.q_RNO_1Z0Z_1\
        );

    \I__6678\ : CascadeMux
    port map (
            O => \N__28201\,
            I => \Lab_UT.didp.Sones_subtractor.q_7_i_1_1_cascade_\
        );

    \I__6677\ : InMux
    port map (
            O => \N__28198\,
            I => \N__28193\
        );

    \I__6676\ : InMux
    port map (
            O => \N__28197\,
            I => \N__28188\
        );

    \I__6675\ : InMux
    port map (
            O => \N__28196\,
            I => \N__28188\
        );

    \I__6674\ : LocalMux
    port map (
            O => \N__28193\,
            I => \N__28185\
        );

    \I__6673\ : LocalMux
    port map (
            O => \N__28188\,
            I => \Lab_UT.didp.Sones_subtractor.q_RNI775L5_1_3\
        );

    \I__6672\ : Odrv4
    port map (
            O => \N__28185\,
            I => \Lab_UT.didp.Sones_subtractor.q_RNI775L5_1_3\
        );

    \I__6671\ : InMux
    port map (
            O => \N__28180\,
            I => \N__28176\
        );

    \I__6670\ : InMux
    port map (
            O => \N__28179\,
            I => \N__28168\
        );

    \I__6669\ : LocalMux
    port map (
            O => \N__28176\,
            I => \N__28165\
        );

    \I__6668\ : CascadeMux
    port map (
            O => \N__28175\,
            I => \N__28162\
        );

    \I__6667\ : InMux
    port map (
            O => \N__28174\,
            I => \N__28156\
        );

    \I__6666\ : InMux
    port map (
            O => \N__28173\,
            I => \N__28156\
        );

    \I__6665\ : InMux
    port map (
            O => \N__28172\,
            I => \N__28151\
        );

    \I__6664\ : InMux
    port map (
            O => \N__28171\,
            I => \N__28151\
        );

    \I__6663\ : LocalMux
    port map (
            O => \N__28168\,
            I => \N__28148\
        );

    \I__6662\ : Span4Mux_v
    port map (
            O => \N__28165\,
            I => \N__28145\
        );

    \I__6661\ : InMux
    port map (
            O => \N__28162\,
            I => \N__28140\
        );

    \I__6660\ : InMux
    port map (
            O => \N__28161\,
            I => \N__28140\
        );

    \I__6659\ : LocalMux
    port map (
            O => \N__28156\,
            I => \Lab_UT.didp.N_82\
        );

    \I__6658\ : LocalMux
    port map (
            O => \N__28151\,
            I => \Lab_UT.didp.N_82\
        );

    \I__6657\ : Odrv4
    port map (
            O => \N__28148\,
            I => \Lab_UT.didp.N_82\
        );

    \I__6656\ : Odrv4
    port map (
            O => \N__28145\,
            I => \Lab_UT.didp.N_82\
        );

    \I__6655\ : LocalMux
    port map (
            O => \N__28140\,
            I => \Lab_UT.didp.N_82\
        );

    \I__6654\ : CascadeMux
    port map (
            O => \N__28129\,
            I => \Lab_UT.didp.Sones_subtractor.un1_q_axb0_cascade_\
        );

    \I__6653\ : InMux
    port map (
            O => \N__28126\,
            I => \N__28120\
        );

    \I__6652\ : InMux
    port map (
            O => \N__28125\,
            I => \N__28117\
        );

    \I__6651\ : InMux
    port map (
            O => \N__28124\,
            I => \N__28112\
        );

    \I__6650\ : InMux
    port map (
            O => \N__28123\,
            I => \N__28112\
        );

    \I__6649\ : LocalMux
    port map (
            O => \N__28120\,
            I => \Lab_UT.didp.Sones_subtractor.N_85\
        );

    \I__6648\ : LocalMux
    port map (
            O => \N__28117\,
            I => \Lab_UT.didp.Sones_subtractor.N_85\
        );

    \I__6647\ : LocalMux
    port map (
            O => \N__28112\,
            I => \Lab_UT.didp.Sones_subtractor.N_85\
        );

    \I__6646\ : InMux
    port map (
            O => \N__28105\,
            I => \N__28099\
        );

    \I__6645\ : InMux
    port map (
            O => \N__28104\,
            I => \N__28096\
        );

    \I__6644\ : CascadeMux
    port map (
            O => \N__28103\,
            I => \N__28093\
        );

    \I__6643\ : CascadeMux
    port map (
            O => \N__28102\,
            I => \N__28089\
        );

    \I__6642\ : LocalMux
    port map (
            O => \N__28099\,
            I => \N__28085\
        );

    \I__6641\ : LocalMux
    port map (
            O => \N__28096\,
            I => \N__28082\
        );

    \I__6640\ : InMux
    port map (
            O => \N__28093\,
            I => \N__28077\
        );

    \I__6639\ : InMux
    port map (
            O => \N__28092\,
            I => \N__28077\
        );

    \I__6638\ : InMux
    port map (
            O => \N__28089\,
            I => \N__28072\
        );

    \I__6637\ : InMux
    port map (
            O => \N__28088\,
            I => \N__28072\
        );

    \I__6636\ : Span4Mux_v
    port map (
            O => \N__28085\,
            I => \N__28067\
        );

    \I__6635\ : Span4Mux_h
    port map (
            O => \N__28082\,
            I => \N__28067\
        );

    \I__6634\ : LocalMux
    port map (
            O => \N__28077\,
            I => \Lab_UT.didp.di_Sones_1\
        );

    \I__6633\ : LocalMux
    port map (
            O => \N__28072\,
            I => \Lab_UT.didp.di_Sones_1\
        );

    \I__6632\ : Odrv4
    port map (
            O => \N__28067\,
            I => \Lab_UT.didp.di_Sones_1\
        );

    \I__6631\ : CascadeMux
    port map (
            O => \N__28060\,
            I => \N__28056\
        );

    \I__6630\ : CascadeMux
    port map (
            O => \N__28059\,
            I => \N__28052\
        );

    \I__6629\ : InMux
    port map (
            O => \N__28056\,
            I => \N__28040\
        );

    \I__6628\ : InMux
    port map (
            O => \N__28055\,
            I => \N__28040\
        );

    \I__6627\ : InMux
    port map (
            O => \N__28052\,
            I => \N__28040\
        );

    \I__6626\ : InMux
    port map (
            O => \N__28051\,
            I => \N__28040\
        );

    \I__6625\ : InMux
    port map (
            O => \N__28050\,
            I => \N__28035\
        );

    \I__6624\ : InMux
    port map (
            O => \N__28049\,
            I => \N__28035\
        );

    \I__6623\ : LocalMux
    port map (
            O => \N__28040\,
            I => \Lab_UT.didp.N_81\
        );

    \I__6622\ : LocalMux
    port map (
            O => \N__28035\,
            I => \Lab_UT.didp.N_81\
        );

    \I__6621\ : InMux
    port map (
            O => \N__28030\,
            I => \N__28027\
        );

    \I__6620\ : LocalMux
    port map (
            O => \N__28027\,
            I => \Lab_UT.didp.Sones_subtractor.un1_q_c2\
        );

    \I__6619\ : InMux
    port map (
            O => \N__28024\,
            I => \N__28016\
        );

    \I__6618\ : InMux
    port map (
            O => \N__28023\,
            I => \N__28013\
        );

    \I__6617\ : CascadeMux
    port map (
            O => \N__28022\,
            I => \N__28010\
        );

    \I__6616\ : CascadeMux
    port map (
            O => \N__28021\,
            I => \N__28007\
        );

    \I__6615\ : InMux
    port map (
            O => \N__28020\,
            I => \N__28002\
        );

    \I__6614\ : InMux
    port map (
            O => \N__28019\,
            I => \N__28002\
        );

    \I__6613\ : LocalMux
    port map (
            O => \N__28016\,
            I => \N__27999\
        );

    \I__6612\ : LocalMux
    port map (
            O => \N__28013\,
            I => \N__27996\
        );

    \I__6611\ : InMux
    port map (
            O => \N__28010\,
            I => \N__27991\
        );

    \I__6610\ : InMux
    port map (
            O => \N__28007\,
            I => \N__27991\
        );

    \I__6609\ : LocalMux
    port map (
            O => \N__28002\,
            I => \Lab_UT.didp.un4_Mtens_ce\
        );

    \I__6608\ : Odrv4
    port map (
            O => \N__27999\,
            I => \Lab_UT.didp.un4_Mtens_ce\
        );

    \I__6607\ : Odrv4
    port map (
            O => \N__27996\,
            I => \Lab_UT.didp.un4_Mtens_ce\
        );

    \I__6606\ : LocalMux
    port map (
            O => \N__27991\,
            I => \Lab_UT.didp.un4_Mtens_ce\
        );

    \I__6605\ : InMux
    port map (
            O => \N__27982\,
            I => \N__27972\
        );

    \I__6604\ : InMux
    port map (
            O => \N__27981\,
            I => \N__27972\
        );

    \I__6603\ : InMux
    port map (
            O => \N__27980\,
            I => \N__27972\
        );

    \I__6602\ : InMux
    port map (
            O => \N__27979\,
            I => \N__27969\
        );

    \I__6601\ : LocalMux
    port map (
            O => \N__27972\,
            I => \Lab_UT.didp.Mtens_subtractor.N_87\
        );

    \I__6600\ : LocalMux
    port map (
            O => \N__27969\,
            I => \Lab_UT.didp.Mtens_subtractor.N_87\
        );

    \I__6599\ : InMux
    port map (
            O => \N__27964\,
            I => \N__27961\
        );

    \I__6598\ : LocalMux
    port map (
            O => \N__27961\,
            I => \Lab_UT.didp.Mtens_subtractor.N_145\
        );

    \I__6597\ : InMux
    port map (
            O => \N__27958\,
            I => \N__27955\
        );

    \I__6596\ : LocalMux
    port map (
            O => \N__27955\,
            I => \N__27952\
        );

    \I__6595\ : Odrv4
    port map (
            O => \N__27952\,
            I => \Lab_UT.didp.Mtens_subtractor.un1_q_c2\
        );

    \I__6594\ : CascadeMux
    port map (
            O => \N__27949\,
            I => \N__27944\
        );

    \I__6593\ : InMux
    port map (
            O => \N__27948\,
            I => \N__27939\
        );

    \I__6592\ : CascadeMux
    port map (
            O => \N__27947\,
            I => \N__27935\
        );

    \I__6591\ : InMux
    port map (
            O => \N__27944\,
            I => \N__27931\
        );

    \I__6590\ : InMux
    port map (
            O => \N__27943\,
            I => \N__27926\
        );

    \I__6589\ : InMux
    port map (
            O => \N__27942\,
            I => \N__27926\
        );

    \I__6588\ : LocalMux
    port map (
            O => \N__27939\,
            I => \N__27923\
        );

    \I__6587\ : InMux
    port map (
            O => \N__27938\,
            I => \N__27920\
        );

    \I__6586\ : InMux
    port map (
            O => \N__27935\,
            I => \N__27917\
        );

    \I__6585\ : InMux
    port map (
            O => \N__27934\,
            I => \N__27914\
        );

    \I__6584\ : LocalMux
    port map (
            O => \N__27931\,
            I => \N__27911\
        );

    \I__6583\ : LocalMux
    port map (
            O => \N__27926\,
            I => \N__27908\
        );

    \I__6582\ : Span4Mux_h
    port map (
            O => \N__27923\,
            I => \N__27905\
        );

    \I__6581\ : LocalMux
    port map (
            O => \N__27920\,
            I => \Lab_UT.didp.di_Mtens_1\
        );

    \I__6580\ : LocalMux
    port map (
            O => \N__27917\,
            I => \Lab_UT.didp.di_Mtens_1\
        );

    \I__6579\ : LocalMux
    port map (
            O => \N__27914\,
            I => \Lab_UT.didp.di_Mtens_1\
        );

    \I__6578\ : Odrv4
    port map (
            O => \N__27911\,
            I => \Lab_UT.didp.di_Mtens_1\
        );

    \I__6577\ : Odrv4
    port map (
            O => \N__27908\,
            I => \Lab_UT.didp.di_Mtens_1\
        );

    \I__6576\ : Odrv4
    port map (
            O => \N__27905\,
            I => \Lab_UT.didp.di_Mtens_1\
        );

    \I__6575\ : CascadeMux
    port map (
            O => \N__27892\,
            I => \Lab_UT.didp.q_RNITOVP_1_cascade_\
        );

    \I__6574\ : IoInMux
    port map (
            O => \N__27889\,
            I => \N__27886\
        );

    \I__6573\ : LocalMux
    port map (
            O => \N__27886\,
            I => \N__27883\
        );

    \I__6572\ : IoSpan4Mux
    port map (
            O => \N__27883\,
            I => \N__27880\
        );

    \I__6571\ : Odrv4
    port map (
            O => \N__27880\,
            I => led_c_1
        );

    \I__6570\ : CascadeMux
    port map (
            O => \N__27877\,
            I => \N__27874\
        );

    \I__6569\ : InMux
    port map (
            O => \N__27874\,
            I => \N__27864\
        );

    \I__6568\ : InMux
    port map (
            O => \N__27873\,
            I => \N__27864\
        );

    \I__6567\ : InMux
    port map (
            O => \N__27872\,
            I => \N__27861\
        );

    \I__6566\ : InMux
    port map (
            O => \N__27871\,
            I => \N__27858\
        );

    \I__6565\ : InMux
    port map (
            O => \N__27870\,
            I => \N__27855\
        );

    \I__6564\ : InMux
    port map (
            O => \N__27869\,
            I => \N__27852\
        );

    \I__6563\ : LocalMux
    port map (
            O => \N__27864\,
            I => \N__27847\
        );

    \I__6562\ : LocalMux
    port map (
            O => \N__27861\,
            I => \N__27847\
        );

    \I__6561\ : LocalMux
    port map (
            O => \N__27858\,
            I => \N__27842\
        );

    \I__6560\ : LocalMux
    port map (
            O => \N__27855\,
            I => \N__27842\
        );

    \I__6559\ : LocalMux
    port map (
            O => \N__27852\,
            I => \N__27837\
        );

    \I__6558\ : Span4Mux_h
    port map (
            O => \N__27847\,
            I => \N__27837\
        );

    \I__6557\ : Odrv12
    port map (
            O => \N__27842\,
            I => \Lab_UT.didp.di_Stens_1\
        );

    \I__6556\ : Odrv4
    port map (
            O => \N__27837\,
            I => \Lab_UT.didp.di_Stens_1\
        );

    \I__6555\ : InMux
    port map (
            O => \N__27832\,
            I => \N__27829\
        );

    \I__6554\ : LocalMux
    port map (
            O => \N__27829\,
            I => \Lab_UT.didp.q_RNI99F11_1\
        );

    \I__6553\ : InMux
    port map (
            O => \N__27826\,
            I => \N__27823\
        );

    \I__6552\ : LocalMux
    port map (
            O => \N__27823\,
            I => \N__27820\
        );

    \I__6551\ : Span4Mux_s3_h
    port map (
            O => \N__27820\,
            I => \N__27817\
        );

    \I__6550\ : Odrv4
    port map (
            O => \N__27817\,
            I => \Lab_UT.dictrl.r_dicLdMtens15\
        );

    \I__6549\ : CascadeMux
    port map (
            O => \N__27814\,
            I => \N__27803\
        );

    \I__6548\ : InMux
    port map (
            O => \N__27813\,
            I => \N__27799\
        );

    \I__6547\ : InMux
    port map (
            O => \N__27812\,
            I => \N__27796\
        );

    \I__6546\ : InMux
    port map (
            O => \N__27811\,
            I => \N__27784\
        );

    \I__6545\ : CascadeMux
    port map (
            O => \N__27810\,
            I => \N__27778\
        );

    \I__6544\ : InMux
    port map (
            O => \N__27809\,
            I => \N__27774\
        );

    \I__6543\ : InMux
    port map (
            O => \N__27808\,
            I => \N__27766\
        );

    \I__6542\ : InMux
    port map (
            O => \N__27807\,
            I => \N__27766\
        );

    \I__6541\ : InMux
    port map (
            O => \N__27806\,
            I => \N__27766\
        );

    \I__6540\ : InMux
    port map (
            O => \N__27803\,
            I => \N__27761\
        );

    \I__6539\ : InMux
    port map (
            O => \N__27802\,
            I => \N__27761\
        );

    \I__6538\ : LocalMux
    port map (
            O => \N__27799\,
            I => \N__27756\
        );

    \I__6537\ : LocalMux
    port map (
            O => \N__27796\,
            I => \N__27756\
        );

    \I__6536\ : InMux
    port map (
            O => \N__27795\,
            I => \N__27749\
        );

    \I__6535\ : InMux
    port map (
            O => \N__27794\,
            I => \N__27749\
        );

    \I__6534\ : InMux
    port map (
            O => \N__27793\,
            I => \N__27749\
        );

    \I__6533\ : InMux
    port map (
            O => \N__27792\,
            I => \N__27740\
        );

    \I__6532\ : InMux
    port map (
            O => \N__27791\,
            I => \N__27740\
        );

    \I__6531\ : InMux
    port map (
            O => \N__27790\,
            I => \N__27735\
        );

    \I__6530\ : InMux
    port map (
            O => \N__27789\,
            I => \N__27735\
        );

    \I__6529\ : CascadeMux
    port map (
            O => \N__27788\,
            I => \N__27732\
        );

    \I__6528\ : InMux
    port map (
            O => \N__27787\,
            I => \N__27726\
        );

    \I__6527\ : LocalMux
    port map (
            O => \N__27784\,
            I => \N__27722\
        );

    \I__6526\ : InMux
    port map (
            O => \N__27783\,
            I => \N__27717\
        );

    \I__6525\ : InMux
    port map (
            O => \N__27782\,
            I => \N__27717\
        );

    \I__6524\ : InMux
    port map (
            O => \N__27781\,
            I => \N__27713\
        );

    \I__6523\ : InMux
    port map (
            O => \N__27778\,
            I => \N__27705\
        );

    \I__6522\ : InMux
    port map (
            O => \N__27777\,
            I => \N__27705\
        );

    \I__6521\ : LocalMux
    port map (
            O => \N__27774\,
            I => \N__27702\
        );

    \I__6520\ : InMux
    port map (
            O => \N__27773\,
            I => \N__27697\
        );

    \I__6519\ : LocalMux
    port map (
            O => \N__27766\,
            I => \N__27692\
        );

    \I__6518\ : LocalMux
    port map (
            O => \N__27761\,
            I => \N__27692\
        );

    \I__6517\ : Span4Mux_v
    port map (
            O => \N__27756\,
            I => \N__27687\
        );

    \I__6516\ : LocalMux
    port map (
            O => \N__27749\,
            I => \N__27687\
        );

    \I__6515\ : InMux
    port map (
            O => \N__27748\,
            I => \N__27684\
        );

    \I__6514\ : InMux
    port map (
            O => \N__27747\,
            I => \N__27677\
        );

    \I__6513\ : InMux
    port map (
            O => \N__27746\,
            I => \N__27677\
        );

    \I__6512\ : InMux
    port map (
            O => \N__27745\,
            I => \N__27677\
        );

    \I__6511\ : LocalMux
    port map (
            O => \N__27740\,
            I => \N__27672\
        );

    \I__6510\ : LocalMux
    port map (
            O => \N__27735\,
            I => \N__27672\
        );

    \I__6509\ : InMux
    port map (
            O => \N__27732\,
            I => \N__27665\
        );

    \I__6508\ : InMux
    port map (
            O => \N__27731\,
            I => \N__27665\
        );

    \I__6507\ : InMux
    port map (
            O => \N__27730\,
            I => \N__27665\
        );

    \I__6506\ : InMux
    port map (
            O => \N__27729\,
            I => \N__27662\
        );

    \I__6505\ : LocalMux
    port map (
            O => \N__27726\,
            I => \N__27659\
        );

    \I__6504\ : InMux
    port map (
            O => \N__27725\,
            I => \N__27656\
        );

    \I__6503\ : Span4Mux_h
    port map (
            O => \N__27722\,
            I => \N__27651\
        );

    \I__6502\ : LocalMux
    port map (
            O => \N__27717\,
            I => \N__27651\
        );

    \I__6501\ : InMux
    port map (
            O => \N__27716\,
            I => \N__27648\
        );

    \I__6500\ : LocalMux
    port map (
            O => \N__27713\,
            I => \N__27640\
        );

    \I__6499\ : InMux
    port map (
            O => \N__27712\,
            I => \N__27637\
        );

    \I__6498\ : InMux
    port map (
            O => \N__27711\,
            I => \N__27632\
        );

    \I__6497\ : InMux
    port map (
            O => \N__27710\,
            I => \N__27632\
        );

    \I__6496\ : LocalMux
    port map (
            O => \N__27705\,
            I => \N__27629\
        );

    \I__6495\ : Span4Mux_h
    port map (
            O => \N__27702\,
            I => \N__27626\
        );

    \I__6494\ : InMux
    port map (
            O => \N__27701\,
            I => \N__27621\
        );

    \I__6493\ : InMux
    port map (
            O => \N__27700\,
            I => \N__27621\
        );

    \I__6492\ : LocalMux
    port map (
            O => \N__27697\,
            I => \N__27612\
        );

    \I__6491\ : Span4Mux_v
    port map (
            O => \N__27692\,
            I => \N__27612\
        );

    \I__6490\ : Span4Mux_h
    port map (
            O => \N__27687\,
            I => \N__27612\
        );

    \I__6489\ : LocalMux
    port map (
            O => \N__27684\,
            I => \N__27612\
        );

    \I__6488\ : LocalMux
    port map (
            O => \N__27677\,
            I => \N__27605\
        );

    \I__6487\ : Span4Mux_h
    port map (
            O => \N__27672\,
            I => \N__27605\
        );

    \I__6486\ : LocalMux
    port map (
            O => \N__27665\,
            I => \N__27605\
        );

    \I__6485\ : LocalMux
    port map (
            O => \N__27662\,
            I => \N__27594\
        );

    \I__6484\ : Span4Mux_h
    port map (
            O => \N__27659\,
            I => \N__27594\
        );

    \I__6483\ : LocalMux
    port map (
            O => \N__27656\,
            I => \N__27594\
        );

    \I__6482\ : Span4Mux_v
    port map (
            O => \N__27651\,
            I => \N__27594\
        );

    \I__6481\ : LocalMux
    port map (
            O => \N__27648\,
            I => \N__27594\
        );

    \I__6480\ : InMux
    port map (
            O => \N__27647\,
            I => \N__27583\
        );

    \I__6479\ : InMux
    port map (
            O => \N__27646\,
            I => \N__27583\
        );

    \I__6478\ : InMux
    port map (
            O => \N__27645\,
            I => \N__27583\
        );

    \I__6477\ : InMux
    port map (
            O => \N__27644\,
            I => \N__27583\
        );

    \I__6476\ : InMux
    port map (
            O => \N__27643\,
            I => \N__27583\
        );

    \I__6475\ : Odrv4
    port map (
            O => \N__27640\,
            I => bu_rx_data_rdy
        );

    \I__6474\ : LocalMux
    port map (
            O => \N__27637\,
            I => bu_rx_data_rdy
        );

    \I__6473\ : LocalMux
    port map (
            O => \N__27632\,
            I => bu_rx_data_rdy
        );

    \I__6472\ : Odrv4
    port map (
            O => \N__27629\,
            I => bu_rx_data_rdy
        );

    \I__6471\ : Odrv4
    port map (
            O => \N__27626\,
            I => bu_rx_data_rdy
        );

    \I__6470\ : LocalMux
    port map (
            O => \N__27621\,
            I => bu_rx_data_rdy
        );

    \I__6469\ : Odrv4
    port map (
            O => \N__27612\,
            I => bu_rx_data_rdy
        );

    \I__6468\ : Odrv4
    port map (
            O => \N__27605\,
            I => bu_rx_data_rdy
        );

    \I__6467\ : Odrv4
    port map (
            O => \N__27594\,
            I => bu_rx_data_rdy
        );

    \I__6466\ : LocalMux
    port map (
            O => \N__27583\,
            I => bu_rx_data_rdy
        );

    \I__6465\ : InMux
    port map (
            O => \N__27562\,
            I => \N__27556\
        );

    \I__6464\ : InMux
    port map (
            O => \N__27561\,
            I => \N__27553\
        );

    \I__6463\ : InMux
    port map (
            O => \N__27560\,
            I => \N__27546\
        );

    \I__6462\ : InMux
    port map (
            O => \N__27559\,
            I => \N__27546\
        );

    \I__6461\ : LocalMux
    port map (
            O => \N__27556\,
            I => \N__27538\
        );

    \I__6460\ : LocalMux
    port map (
            O => \N__27553\,
            I => \N__27535\
        );

    \I__6459\ : InMux
    port map (
            O => \N__27552\,
            I => \N__27532\
        );

    \I__6458\ : InMux
    port map (
            O => \N__27551\,
            I => \N__27529\
        );

    \I__6457\ : LocalMux
    port map (
            O => \N__27546\,
            I => \N__27526\
        );

    \I__6456\ : InMux
    port map (
            O => \N__27545\,
            I => \N__27521\
        );

    \I__6455\ : InMux
    port map (
            O => \N__27544\,
            I => \N__27521\
        );

    \I__6454\ : InMux
    port map (
            O => \N__27543\,
            I => \N__27518\
        );

    \I__6453\ : InMux
    port map (
            O => \N__27542\,
            I => \N__27512\
        );

    \I__6452\ : InMux
    port map (
            O => \N__27541\,
            I => \N__27512\
        );

    \I__6451\ : Span4Mux_v
    port map (
            O => \N__27538\,
            I => \N__27507\
        );

    \I__6450\ : Span4Mux_v
    port map (
            O => \N__27535\,
            I => \N__27504\
        );

    \I__6449\ : LocalMux
    port map (
            O => \N__27532\,
            I => \N__27501\
        );

    \I__6448\ : LocalMux
    port map (
            O => \N__27529\,
            I => \N__27498\
        );

    \I__6447\ : Span4Mux_v
    port map (
            O => \N__27526\,
            I => \N__27493\
        );

    \I__6446\ : LocalMux
    port map (
            O => \N__27521\,
            I => \N__27493\
        );

    \I__6445\ : LocalMux
    port map (
            O => \N__27518\,
            I => \N__27490\
        );

    \I__6444\ : InMux
    port map (
            O => \N__27517\,
            I => \N__27487\
        );

    \I__6443\ : LocalMux
    port map (
            O => \N__27512\,
            I => \N__27484\
        );

    \I__6442\ : CascadeMux
    port map (
            O => \N__27511\,
            I => \N__27479\
        );

    \I__6441\ : CascadeMux
    port map (
            O => \N__27510\,
            I => \N__27476\
        );

    \I__6440\ : Span4Mux_h
    port map (
            O => \N__27507\,
            I => \N__27468\
        );

    \I__6439\ : Span4Mux_s2_h
    port map (
            O => \N__27504\,
            I => \N__27468\
        );

    \I__6438\ : Span4Mux_v
    port map (
            O => \N__27501\,
            I => \N__27468\
        );

    \I__6437\ : Span4Mux_v
    port map (
            O => \N__27498\,
            I => \N__27461\
        );

    \I__6436\ : Span4Mux_h
    port map (
            O => \N__27493\,
            I => \N__27461\
        );

    \I__6435\ : Span4Mux_s3_h
    port map (
            O => \N__27490\,
            I => \N__27461\
        );

    \I__6434\ : LocalMux
    port map (
            O => \N__27487\,
            I => \N__27456\
        );

    \I__6433\ : Span4Mux_s3_h
    port map (
            O => \N__27484\,
            I => \N__27456\
        );

    \I__6432\ : InMux
    port map (
            O => \N__27483\,
            I => \N__27445\
        );

    \I__6431\ : InMux
    port map (
            O => \N__27482\,
            I => \N__27445\
        );

    \I__6430\ : InMux
    port map (
            O => \N__27479\,
            I => \N__27445\
        );

    \I__6429\ : InMux
    port map (
            O => \N__27476\,
            I => \N__27445\
        );

    \I__6428\ : InMux
    port map (
            O => \N__27475\,
            I => \N__27445\
        );

    \I__6427\ : Odrv4
    port map (
            O => \N__27468\,
            I => \Lab_UT.dictrl.de_num_0\
        );

    \I__6426\ : Odrv4
    port map (
            O => \N__27461\,
            I => \Lab_UT.dictrl.de_num_0\
        );

    \I__6425\ : Odrv4
    port map (
            O => \N__27456\,
            I => \Lab_UT.dictrl.de_num_0\
        );

    \I__6424\ : LocalMux
    port map (
            O => \N__27445\,
            I => \Lab_UT.dictrl.de_num_0\
        );

    \I__6423\ : InMux
    port map (
            O => \N__27436\,
            I => \N__27430\
        );

    \I__6422\ : InMux
    port map (
            O => \N__27435\,
            I => \N__27430\
        );

    \I__6421\ : LocalMux
    port map (
            O => \N__27430\,
            I => \N__27427\
        );

    \I__6420\ : Odrv4
    port map (
            O => \N__27427\,
            I => \Lab_UT.dicLdMones_latmux\
        );

    \I__6419\ : InMux
    port map (
            O => \N__27424\,
            I => \N__27421\
        );

    \I__6418\ : LocalMux
    port map (
            O => \N__27421\,
            I => \N__27418\
        );

    \I__6417\ : Odrv12
    port map (
            O => \N__27418\,
            I => \Lab_UT.displayAlarmZ0Z_6\
        );

    \I__6416\ : InMux
    port map (
            O => \N__27415\,
            I => \N__27408\
        );

    \I__6415\ : InMux
    port map (
            O => \N__27414\,
            I => \N__27408\
        );

    \I__6414\ : InMux
    port map (
            O => \N__27413\,
            I => \N__27405\
        );

    \I__6413\ : LocalMux
    port map (
            O => \N__27408\,
            I => \N__27402\
        );

    \I__6412\ : LocalMux
    port map (
            O => \N__27405\,
            I => \N__27399\
        );

    \I__6411\ : Span4Mux_s3_h
    port map (
            O => \N__27402\,
            I => \N__27396\
        );

    \I__6410\ : Span4Mux_s2_h
    port map (
            O => \N__27399\,
            I => \N__27392\
        );

    \I__6409\ : Span4Mux_v
    port map (
            O => \N__27396\,
            I => \N__27389\
        );

    \I__6408\ : CascadeMux
    port map (
            O => \N__27395\,
            I => \N__27385\
        );

    \I__6407\ : Span4Mux_v
    port map (
            O => \N__27392\,
            I => \N__27382\
        );

    \I__6406\ : Sp12to4
    port map (
            O => \N__27389\,
            I => \N__27379\
        );

    \I__6405\ : InMux
    port map (
            O => \N__27388\,
            I => \N__27374\
        );

    \I__6404\ : InMux
    port map (
            O => \N__27385\,
            I => \N__27374\
        );

    \I__6403\ : Odrv4
    port map (
            O => \N__27382\,
            I => \Lab_UT.alarm_armed\
        );

    \I__6402\ : Odrv12
    port map (
            O => \N__27379\,
            I => \Lab_UT.alarm_armed\
        );

    \I__6401\ : LocalMux
    port map (
            O => \N__27374\,
            I => \Lab_UT.alarm_armed\
        );

    \I__6400\ : InMux
    port map (
            O => \N__27367\,
            I => \N__27364\
        );

    \I__6399\ : LocalMux
    port map (
            O => \N__27364\,
            I => \N__27361\
        );

    \I__6398\ : Span4Mux_v
    port map (
            O => \N__27361\,
            I => \N__27358\
        );

    \I__6397\ : Odrv4
    port map (
            O => \N__27358\,
            I => \Lab_UT.displayAlarmZ0Z_4\
        );

    \I__6396\ : InMux
    port map (
            O => \N__27355\,
            I => \N__27346\
        );

    \I__6395\ : InMux
    port map (
            O => \N__27354\,
            I => \N__27346\
        );

    \I__6394\ : InMux
    port map (
            O => \N__27353\,
            I => \N__27346\
        );

    \I__6393\ : LocalMux
    port map (
            O => \N__27346\,
            I => \N__27342\
        );

    \I__6392\ : InMux
    port map (
            O => \N__27345\,
            I => \N__27338\
        );

    \I__6391\ : Span4Mux_h
    port map (
            O => \N__27342\,
            I => \N__27335\
        );

    \I__6390\ : InMux
    port map (
            O => \N__27341\,
            I => \N__27332\
        );

    \I__6389\ : LocalMux
    port map (
            O => \N__27338\,
            I => \Lab_UT.alarm_match\
        );

    \I__6388\ : Odrv4
    port map (
            O => \N__27335\,
            I => \Lab_UT.alarm_match\
        );

    \I__6387\ : LocalMux
    port map (
            O => \N__27332\,
            I => \Lab_UT.alarm_match\
        );

    \I__6386\ : CascadeMux
    port map (
            O => \N__27325\,
            I => \N__27321\
        );

    \I__6385\ : InMux
    port map (
            O => \N__27324\,
            I => \N__27316\
        );

    \I__6384\ : InMux
    port map (
            O => \N__27321\,
            I => \N__27316\
        );

    \I__6383\ : LocalMux
    port map (
            O => \N__27316\,
            I => \Lab_UT.dicLdMones\
        );

    \I__6382\ : InMux
    port map (
            O => \N__27313\,
            I => \N__27310\
        );

    \I__6381\ : LocalMux
    port map (
            O => \N__27310\,
            I => \N__27307\
        );

    \I__6380\ : Span4Mux_h
    port map (
            O => \N__27307\,
            I => \N__27304\
        );

    \I__6379\ : Odrv4
    port map (
            O => \N__27304\,
            I => \Lab_UT.dictrl.r_dicLdMtens14\
        );

    \I__6378\ : InMux
    port map (
            O => \N__27301\,
            I => \N__27289\
        );

    \I__6377\ : InMux
    port map (
            O => \N__27300\,
            I => \N__27286\
        );

    \I__6376\ : InMux
    port map (
            O => \N__27299\,
            I => \N__27281\
        );

    \I__6375\ : InMux
    port map (
            O => \N__27298\,
            I => \N__27278\
        );

    \I__6374\ : InMux
    port map (
            O => \N__27297\,
            I => \N__27271\
        );

    \I__6373\ : InMux
    port map (
            O => \N__27296\,
            I => \N__27271\
        );

    \I__6372\ : InMux
    port map (
            O => \N__27295\,
            I => \N__27264\
        );

    \I__6371\ : InMux
    port map (
            O => \N__27294\,
            I => \N__27264\
        );

    \I__6370\ : InMux
    port map (
            O => \N__27293\,
            I => \N__27264\
        );

    \I__6369\ : InMux
    port map (
            O => \N__27292\,
            I => \N__27261\
        );

    \I__6368\ : LocalMux
    port map (
            O => \N__27289\,
            I => \N__27258\
        );

    \I__6367\ : LocalMux
    port map (
            O => \N__27286\,
            I => \N__27255\
        );

    \I__6366\ : InMux
    port map (
            O => \N__27285\,
            I => \N__27250\
        );

    \I__6365\ : InMux
    port map (
            O => \N__27284\,
            I => \N__27250\
        );

    \I__6364\ : LocalMux
    port map (
            O => \N__27281\,
            I => \N__27243\
        );

    \I__6363\ : LocalMux
    port map (
            O => \N__27278\,
            I => \N__27240\
        );

    \I__6362\ : InMux
    port map (
            O => \N__27277\,
            I => \N__27235\
        );

    \I__6361\ : InMux
    port map (
            O => \N__27276\,
            I => \N__27235\
        );

    \I__6360\ : LocalMux
    port map (
            O => \N__27271\,
            I => \N__27232\
        );

    \I__6359\ : LocalMux
    port map (
            O => \N__27264\,
            I => \N__27227\
        );

    \I__6358\ : LocalMux
    port map (
            O => \N__27261\,
            I => \N__27227\
        );

    \I__6357\ : Span4Mux_h
    port map (
            O => \N__27258\,
            I => \N__27220\
        );

    \I__6356\ : Span4Mux_v
    port map (
            O => \N__27255\,
            I => \N__27220\
        );

    \I__6355\ : LocalMux
    port map (
            O => \N__27250\,
            I => \N__27220\
        );

    \I__6354\ : InMux
    port map (
            O => \N__27249\,
            I => \N__27213\
        );

    \I__6353\ : InMux
    port map (
            O => \N__27248\,
            I => \N__27213\
        );

    \I__6352\ : InMux
    port map (
            O => \N__27247\,
            I => \N__27213\
        );

    \I__6351\ : InMux
    port map (
            O => \N__27246\,
            I => \N__27206\
        );

    \I__6350\ : Span4Mux_h
    port map (
            O => \N__27243\,
            I => \N__27201\
        );

    \I__6349\ : Span4Mux_s3_h
    port map (
            O => \N__27240\,
            I => \N__27201\
        );

    \I__6348\ : LocalMux
    port map (
            O => \N__27235\,
            I => \N__27194\
        );

    \I__6347\ : Span4Mux_s3_h
    port map (
            O => \N__27232\,
            I => \N__27194\
        );

    \I__6346\ : Span4Mux_h
    port map (
            O => \N__27227\,
            I => \N__27194\
        );

    \I__6345\ : Span4Mux_h
    port map (
            O => \N__27220\,
            I => \N__27189\
        );

    \I__6344\ : LocalMux
    port map (
            O => \N__27213\,
            I => \N__27189\
        );

    \I__6343\ : InMux
    port map (
            O => \N__27212\,
            I => \N__27180\
        );

    \I__6342\ : InMux
    port map (
            O => \N__27211\,
            I => \N__27180\
        );

    \I__6341\ : InMux
    port map (
            O => \N__27210\,
            I => \N__27180\
        );

    \I__6340\ : InMux
    port map (
            O => \N__27209\,
            I => \N__27180\
        );

    \I__6339\ : LocalMux
    port map (
            O => \N__27206\,
            I => \Lab_UT.dictrl.de_num0to5_1\
        );

    \I__6338\ : Odrv4
    port map (
            O => \N__27201\,
            I => \Lab_UT.dictrl.de_num0to5_1\
        );

    \I__6337\ : Odrv4
    port map (
            O => \N__27194\,
            I => \Lab_UT.dictrl.de_num0to5_1\
        );

    \I__6336\ : Odrv4
    port map (
            O => \N__27189\,
            I => \Lab_UT.dictrl.de_num0to5_1\
        );

    \I__6335\ : LocalMux
    port map (
            O => \N__27180\,
            I => \Lab_UT.dictrl.de_num0to5_1\
        );

    \I__6334\ : CascadeMux
    port map (
            O => \N__27169\,
            I => \Lab_UT.dicLdMtens_latmux_cascade_\
        );

    \I__6333\ : InMux
    port map (
            O => \N__27166\,
            I => \N__27163\
        );

    \I__6332\ : LocalMux
    port map (
            O => \N__27163\,
            I => \N__27156\
        );

    \I__6331\ : InMux
    port map (
            O => \N__27162\,
            I => \N__27153\
        );

    \I__6330\ : InMux
    port map (
            O => \N__27161\,
            I => \N__27148\
        );

    \I__6329\ : InMux
    port map (
            O => \N__27160\,
            I => \N__27148\
        );

    \I__6328\ : InMux
    port map (
            O => \N__27159\,
            I => \N__27145\
        );

    \I__6327\ : Span4Mux_s2_h
    port map (
            O => \N__27156\,
            I => \N__27142\
        );

    \I__6326\ : LocalMux
    port map (
            O => \N__27153\,
            I => \N__27139\
        );

    \I__6325\ : LocalMux
    port map (
            O => \N__27148\,
            I => \Lab_UT.didp.di_Stens_2\
        );

    \I__6324\ : LocalMux
    port map (
            O => \N__27145\,
            I => \Lab_UT.didp.di_Stens_2\
        );

    \I__6323\ : Odrv4
    port map (
            O => \N__27142\,
            I => \Lab_UT.didp.di_Stens_2\
        );

    \I__6322\ : Odrv4
    port map (
            O => \N__27139\,
            I => \Lab_UT.didp.di_Stens_2\
        );

    \I__6321\ : CascadeMux
    port map (
            O => \N__27130\,
            I => \N__27127\
        );

    \I__6320\ : InMux
    port map (
            O => \N__27127\,
            I => \N__27123\
        );

    \I__6319\ : InMux
    port map (
            O => \N__27126\,
            I => \N__27120\
        );

    \I__6318\ : LocalMux
    port map (
            O => \N__27123\,
            I => \N__27115\
        );

    \I__6317\ : LocalMux
    port map (
            O => \N__27120\,
            I => \N__27112\
        );

    \I__6316\ : InMux
    port map (
            O => \N__27119\,
            I => \N__27109\
        );

    \I__6315\ : InMux
    port map (
            O => \N__27118\,
            I => \N__27106\
        );

    \I__6314\ : Span4Mux_s2_h
    port map (
            O => \N__27115\,
            I => \N__27103\
        );

    \I__6313\ : Span4Mux_h
    port map (
            O => \N__27112\,
            I => \N__27100\
        );

    \I__6312\ : LocalMux
    port map (
            O => \N__27109\,
            I => \Lab_UT.didp.di_Stens_3\
        );

    \I__6311\ : LocalMux
    port map (
            O => \N__27106\,
            I => \Lab_UT.didp.di_Stens_3\
        );

    \I__6310\ : Odrv4
    port map (
            O => \N__27103\,
            I => \Lab_UT.didp.di_Stens_3\
        );

    \I__6309\ : Odrv4
    port map (
            O => \N__27100\,
            I => \Lab_UT.didp.di_Stens_3\
        );

    \I__6308\ : CascadeMux
    port map (
            O => \N__27091\,
            I => \N__27086\
        );

    \I__6307\ : CascadeMux
    port map (
            O => \N__27090\,
            I => \N__27082\
        );

    \I__6306\ : CascadeMux
    port map (
            O => \N__27089\,
            I => \N__27078\
        );

    \I__6305\ : InMux
    port map (
            O => \N__27086\,
            I => \N__27075\
        );

    \I__6304\ : InMux
    port map (
            O => \N__27085\,
            I => \N__27068\
        );

    \I__6303\ : InMux
    port map (
            O => \N__27082\,
            I => \N__27068\
        );

    \I__6302\ : InMux
    port map (
            O => \N__27081\,
            I => \N__27068\
        );

    \I__6301\ : InMux
    port map (
            O => \N__27078\,
            I => \N__27065\
        );

    \I__6300\ : LocalMux
    port map (
            O => \N__27075\,
            I => \N__27062\
        );

    \I__6299\ : LocalMux
    port map (
            O => \N__27068\,
            I => \N__27059\
        );

    \I__6298\ : LocalMux
    port map (
            O => \N__27065\,
            I => \Lab_UT.didp.un6_Mtens_ce\
        );

    \I__6297\ : Odrv12
    port map (
            O => \N__27062\,
            I => \Lab_UT.didp.un6_Mtens_ce\
        );

    \I__6296\ : Odrv4
    port map (
            O => \N__27059\,
            I => \Lab_UT.didp.un6_Mtens_ce\
        );

    \I__6295\ : InMux
    port map (
            O => \N__27052\,
            I => \N__27047\
        );

    \I__6294\ : InMux
    port map (
            O => \N__27051\,
            I => \N__27040\
        );

    \I__6293\ : InMux
    port map (
            O => \N__27050\,
            I => \N__27037\
        );

    \I__6292\ : LocalMux
    port map (
            O => \N__27047\,
            I => \N__27034\
        );

    \I__6291\ : InMux
    port map (
            O => \N__27046\,
            I => \N__27025\
        );

    \I__6290\ : InMux
    port map (
            O => \N__27045\,
            I => \N__27025\
        );

    \I__6289\ : InMux
    port map (
            O => \N__27044\,
            I => \N__27025\
        );

    \I__6288\ : InMux
    port map (
            O => \N__27043\,
            I => \N__27025\
        );

    \I__6287\ : LocalMux
    port map (
            O => \N__27040\,
            I => \Lab_UT.didp.un3_Mtens_rst\
        );

    \I__6286\ : LocalMux
    port map (
            O => \N__27037\,
            I => \Lab_UT.didp.un3_Mtens_rst\
        );

    \I__6285\ : Odrv4
    port map (
            O => \N__27034\,
            I => \Lab_UT.didp.un3_Mtens_rst\
        );

    \I__6284\ : LocalMux
    port map (
            O => \N__27025\,
            I => \Lab_UT.didp.un3_Mtens_rst\
        );

    \I__6283\ : InMux
    port map (
            O => \N__27016\,
            I => \N__27013\
        );

    \I__6282\ : LocalMux
    port map (
            O => \N__27013\,
            I => \N__27010\
        );

    \I__6281\ : Odrv4
    port map (
            O => \N__27010\,
            I => \Lab_UT.didp.Mtens_subtractor.q_RNO_2Z0Z_1\
        );

    \I__6280\ : CascadeMux
    port map (
            O => \N__27007\,
            I => \N__27003\
        );

    \I__6279\ : InMux
    port map (
            O => \N__27006\,
            I => \N__26995\
        );

    \I__6278\ : InMux
    port map (
            O => \N__27003\,
            I => \N__26995\
        );

    \I__6277\ : InMux
    port map (
            O => \N__27002\,
            I => \N__26995\
        );

    \I__6276\ : LocalMux
    port map (
            O => \N__26995\,
            I => \Lab_UT.dicLdMtens\
        );

    \I__6275\ : CascadeMux
    port map (
            O => \N__26992\,
            I => \N__26989\
        );

    \I__6274\ : InMux
    port map (
            O => \N__26989\,
            I => \N__26983\
        );

    \I__6273\ : InMux
    port map (
            O => \N__26988\,
            I => \N__26983\
        );

    \I__6272\ : LocalMux
    port map (
            O => \N__26983\,
            I => \Lab_UT.dicLdMtens_latmux\
        );

    \I__6271\ : InMux
    port map (
            O => \N__26980\,
            I => \N__26977\
        );

    \I__6270\ : LocalMux
    port map (
            O => \N__26977\,
            I => \Lab_UT.didp.Mtens_subtractor.N_147\
        );

    \I__6269\ : CascadeMux
    port map (
            O => \N__26974\,
            I => \Lab_UT.didp.Mtens_subtractor.q_RNO_0_3_2_cascade_\
        );

    \I__6268\ : InMux
    port map (
            O => \N__26971\,
            I => \N__26962\
        );

    \I__6267\ : InMux
    port map (
            O => \N__26970\,
            I => \N__26962\
        );

    \I__6266\ : InMux
    port map (
            O => \N__26969\,
            I => \N__26962\
        );

    \I__6265\ : LocalMux
    port map (
            O => \N__26962\,
            I => \N__26957\
        );

    \I__6264\ : InMux
    port map (
            O => \N__26961\,
            I => \N__26954\
        );

    \I__6263\ : CascadeMux
    port map (
            O => \N__26960\,
            I => \N__26951\
        );

    \I__6262\ : Span4Mux_h
    port map (
            O => \N__26957\,
            I => \N__26947\
        );

    \I__6261\ : LocalMux
    port map (
            O => \N__26954\,
            I => \N__26944\
        );

    \I__6260\ : InMux
    port map (
            O => \N__26951\,
            I => \N__26939\
        );

    \I__6259\ : InMux
    port map (
            O => \N__26950\,
            I => \N__26939\
        );

    \I__6258\ : Odrv4
    port map (
            O => \N__26947\,
            I => \Lab_UT.didp.N_83\
        );

    \I__6257\ : Odrv4
    port map (
            O => \N__26944\,
            I => \Lab_UT.didp.N_83\
        );

    \I__6256\ : LocalMux
    port map (
            O => \N__26939\,
            I => \Lab_UT.didp.N_83\
        );

    \I__6255\ : CascadeMux
    port map (
            O => \N__26932\,
            I => \Lab_UT.didp.un3_Mtens_rst_cascade_\
        );

    \I__6254\ : InMux
    port map (
            O => \N__26929\,
            I => \N__26926\
        );

    \I__6253\ : LocalMux
    port map (
            O => \N__26926\,
            I => \N__26923\
        );

    \I__6252\ : Span4Mux_v
    port map (
            O => \N__26923\,
            I => \N__26920\
        );

    \I__6251\ : Span4Mux_h
    port map (
            O => \N__26920\,
            I => \N__26915\
        );

    \I__6250\ : InMux
    port map (
            O => \N__26919\,
            I => \N__26910\
        );

    \I__6249\ : InMux
    port map (
            O => \N__26918\,
            I => \N__26910\
        );

    \I__6248\ : Span4Mux_h
    port map (
            O => \N__26915\,
            I => \N__26907\
        );

    \I__6247\ : LocalMux
    port map (
            O => \N__26910\,
            I => \Lab_UT.didp.q_RNI775L5_3\
        );

    \I__6246\ : Odrv4
    port map (
            O => \N__26907\,
            I => \Lab_UT.didp.q_RNI775L5_3\
        );

    \I__6245\ : CascadeMux
    port map (
            O => \N__26902\,
            I => \Lab_UT.didp.Mtens_subtractor.un1_q_axb0_cascade_\
        );

    \I__6244\ : CascadeMux
    port map (
            O => \N__26899\,
            I => \N__26896\
        );

    \I__6243\ : InMux
    port map (
            O => \N__26896\,
            I => \N__26893\
        );

    \I__6242\ : LocalMux
    port map (
            O => \N__26893\,
            I => \Lab_UT.didp.Mtens_ce\
        );

    \I__6241\ : CascadeMux
    port map (
            O => \N__26890\,
            I => \N__26887\
        );

    \I__6240\ : InMux
    port map (
            O => \N__26887\,
            I => \N__26883\
        );

    \I__6239\ : InMux
    port map (
            O => \N__26886\,
            I => \N__26880\
        );

    \I__6238\ : LocalMux
    port map (
            O => \N__26883\,
            I => \N__26877\
        );

    \I__6237\ : LocalMux
    port map (
            O => \N__26880\,
            I => \N__26874\
        );

    \I__6236\ : Span4Mux_v
    port map (
            O => \N__26877\,
            I => \N__26867\
        );

    \I__6235\ : Span4Mux_v
    port map (
            O => \N__26874\,
            I => \N__26864\
        );

    \I__6234\ : InMux
    port map (
            O => \N__26873\,
            I => \N__26861\
        );

    \I__6233\ : InMux
    port map (
            O => \N__26872\,
            I => \N__26854\
        );

    \I__6232\ : InMux
    port map (
            O => \N__26871\,
            I => \N__26854\
        );

    \I__6231\ : InMux
    port map (
            O => \N__26870\,
            I => \N__26854\
        );

    \I__6230\ : Span4Mux_h
    port map (
            O => \N__26867\,
            I => \N__26851\
        );

    \I__6229\ : Sp12to4
    port map (
            O => \N__26864\,
            I => \N__26846\
        );

    \I__6228\ : LocalMux
    port map (
            O => \N__26861\,
            I => \N__26846\
        );

    \I__6227\ : LocalMux
    port map (
            O => \N__26854\,
            I => \Lab_UT.di_Mtens_2\
        );

    \I__6226\ : Odrv4
    port map (
            O => \N__26851\,
            I => \Lab_UT.di_Mtens_2\
        );

    \I__6225\ : Odrv12
    port map (
            O => \N__26846\,
            I => \Lab_UT.di_Mtens_2\
        );

    \I__6224\ : CascadeMux
    port map (
            O => \N__26839\,
            I => \Lab_UT.didp.Mtens_ce_cascade_\
        );

    \I__6223\ : CascadeMux
    port map (
            O => \N__26836\,
            I => \Lab_UT.didp.Mtens_subtractor.q_RNO_0_2_3_cascade_\
        );

    \I__6222\ : InMux
    port map (
            O => \N__26833\,
            I => \N__26828\
        );

    \I__6221\ : InMux
    port map (
            O => \N__26832\,
            I => \N__26825\
        );

    \I__6220\ : CascadeMux
    port map (
            O => \N__26831\,
            I => \N__26821\
        );

    \I__6219\ : LocalMux
    port map (
            O => \N__26828\,
            I => \N__26818\
        );

    \I__6218\ : LocalMux
    port map (
            O => \N__26825\,
            I => \N__26815\
        );

    \I__6217\ : InMux
    port map (
            O => \N__26824\,
            I => \N__26810\
        );

    \I__6216\ : InMux
    port map (
            O => \N__26821\,
            I => \N__26810\
        );

    \I__6215\ : Span4Mux_h
    port map (
            O => \N__26818\,
            I => \N__26807\
        );

    \I__6214\ : Odrv12
    port map (
            O => \N__26815\,
            I => \Lab_UT.didp.di_Mtens_3\
        );

    \I__6213\ : LocalMux
    port map (
            O => \N__26810\,
            I => \Lab_UT.didp.di_Mtens_3\
        );

    \I__6212\ : Odrv4
    port map (
            O => \N__26807\,
            I => \Lab_UT.didp.di_Mtens_3\
        );

    \I__6211\ : InMux
    port map (
            O => \N__26800\,
            I => \N__26797\
        );

    \I__6210\ : LocalMux
    port map (
            O => \N__26797\,
            I => \N__26791\
        );

    \I__6209\ : InMux
    port map (
            O => \N__26796\,
            I => \N__26786\
        );

    \I__6208\ : InMux
    port map (
            O => \N__26795\,
            I => \N__26786\
        );

    \I__6207\ : InMux
    port map (
            O => \N__26794\,
            I => \N__26781\
        );

    \I__6206\ : Span4Mux_h
    port map (
            O => \N__26791\,
            I => \N__26778\
        );

    \I__6205\ : LocalMux
    port map (
            O => \N__26786\,
            I => \N__26775\
        );

    \I__6204\ : InMux
    port map (
            O => \N__26785\,
            I => \N__26770\
        );

    \I__6203\ : InMux
    port map (
            O => \N__26784\,
            I => \N__26770\
        );

    \I__6202\ : LocalMux
    port map (
            O => \N__26781\,
            I => \o_One_Sec_Pulse\
        );

    \I__6201\ : Odrv4
    port map (
            O => \N__26778\,
            I => \o_One_Sec_Pulse\
        );

    \I__6200\ : Odrv12
    port map (
            O => \N__26775\,
            I => \o_One_Sec_Pulse\
        );

    \I__6199\ : LocalMux
    port map (
            O => \N__26770\,
            I => \o_One_Sec_Pulse\
        );

    \I__6198\ : InMux
    port map (
            O => \N__26761\,
            I => \N__26757\
        );

    \I__6197\ : InMux
    port map (
            O => \N__26760\,
            I => \N__26754\
        );

    \I__6196\ : LocalMux
    port map (
            O => \N__26757\,
            I => \N__26749\
        );

    \I__6195\ : LocalMux
    port map (
            O => \N__26754\,
            I => \N__26749\
        );

    \I__6194\ : Span4Mux_s3_h
    port map (
            O => \N__26749\,
            I => \N__26745\
        );

    \I__6193\ : InMux
    port map (
            O => \N__26748\,
            I => \N__26742\
        );

    \I__6192\ : Span4Mux_h
    port map (
            O => \N__26745\,
            I => \N__26739\
        );

    \I__6191\ : LocalMux
    port map (
            O => \N__26742\,
            I => \uu0_sec_clkD\
        );

    \I__6190\ : Odrv4
    port map (
            O => \N__26739\,
            I => \uu0_sec_clkD\
        );

    \I__6189\ : InMux
    port map (
            O => \N__26734\,
            I => \N__26726\
        );

    \I__6188\ : InMux
    port map (
            O => \N__26733\,
            I => \N__26719\
        );

    \I__6187\ : InMux
    port map (
            O => \N__26732\,
            I => \N__26719\
        );

    \I__6186\ : InMux
    port map (
            O => \N__26731\,
            I => \N__26719\
        );

    \I__6185\ : InMux
    port map (
            O => \N__26730\,
            I => \N__26714\
        );

    \I__6184\ : InMux
    port map (
            O => \N__26729\,
            I => \N__26714\
        );

    \I__6183\ : LocalMux
    port map (
            O => \N__26726\,
            I => \N__26710\
        );

    \I__6182\ : LocalMux
    port map (
            O => \N__26719\,
            I => \N__26705\
        );

    \I__6181\ : LocalMux
    port map (
            O => \N__26714\,
            I => \N__26705\
        );

    \I__6180\ : InMux
    port map (
            O => \N__26713\,
            I => \N__26702\
        );

    \I__6179\ : Span4Mux_h
    port map (
            O => \N__26710\,
            I => \N__26699\
        );

    \I__6178\ : Span4Mux_v
    port map (
            O => \N__26705\,
            I => \N__26696\
        );

    \I__6177\ : LocalMux
    port map (
            O => \N__26702\,
            I => \N__26693\
        );

    \I__6176\ : Span4Mux_v
    port map (
            O => \N__26699\,
            I => \N__26688\
        );

    \I__6175\ : Span4Mux_h
    port map (
            O => \N__26696\,
            I => \N__26688\
        );

    \I__6174\ : Span12Mux_s8_h
    port map (
            O => \N__26693\,
            I => \N__26685\
        );

    \I__6173\ : Odrv4
    port map (
            O => \N__26688\,
            I => \oneSecStrb\
        );

    \I__6172\ : Odrv12
    port map (
            O => \N__26685\,
            I => \oneSecStrb\
        );

    \I__6171\ : InMux
    port map (
            O => \N__26680\,
            I => \N__26668\
        );

    \I__6170\ : InMux
    port map (
            O => \N__26679\,
            I => \N__26668\
        );

    \I__6169\ : InMux
    port map (
            O => \N__26678\,
            I => \N__26668\
        );

    \I__6168\ : InMux
    port map (
            O => \N__26677\,
            I => \N__26662\
        );

    \I__6167\ : InMux
    port map (
            O => \N__26676\,
            I => \N__26662\
        );

    \I__6166\ : InMux
    port map (
            O => \N__26675\,
            I => \N__26659\
        );

    \I__6165\ : LocalMux
    port map (
            O => \N__26668\,
            I => \N__26656\
        );

    \I__6164\ : InMux
    port map (
            O => \N__26667\,
            I => \N__26653\
        );

    \I__6163\ : LocalMux
    port map (
            O => \N__26662\,
            I => \N__26646\
        );

    \I__6162\ : LocalMux
    port map (
            O => \N__26659\,
            I => \N__26646\
        );

    \I__6161\ : Span4Mux_s3_h
    port map (
            O => \N__26656\,
            I => \N__26646\
        );

    \I__6160\ : LocalMux
    port map (
            O => \N__26653\,
            I => \Lab_UT.ld_enable_dicRun\
        );

    \I__6159\ : Odrv4
    port map (
            O => \N__26646\,
            I => \Lab_UT.ld_enable_dicRun\
        );

    \I__6158\ : CascadeMux
    port map (
            O => \N__26641\,
            I => \Lab_UT.didp.N_84_cascade_\
        );

    \I__6157\ : InMux
    port map (
            O => \N__26638\,
            I => \N__26631\
        );

    \I__6156\ : InMux
    port map (
            O => \N__26637\,
            I => \N__26631\
        );

    \I__6155\ : InMux
    port map (
            O => \N__26636\,
            I => \N__26628\
        );

    \I__6154\ : LocalMux
    port map (
            O => \N__26631\,
            I => \Lab_UT.didp.Sones_subtractor.un8_Mtens_ce\
        );

    \I__6153\ : LocalMux
    port map (
            O => \N__26628\,
            I => \Lab_UT.didp.Sones_subtractor.un8_Mtens_ce\
        );

    \I__6152\ : InMux
    port map (
            O => \N__26623\,
            I => \N__26611\
        );

    \I__6151\ : InMux
    port map (
            O => \N__26622\,
            I => \N__26611\
        );

    \I__6150\ : InMux
    port map (
            O => \N__26621\,
            I => \N__26611\
        );

    \I__6149\ : InMux
    port map (
            O => \N__26620\,
            I => \N__26611\
        );

    \I__6148\ : LocalMux
    port map (
            O => \N__26611\,
            I => \N__26608\
        );

    \I__6147\ : Odrv4
    port map (
            O => \N__26608\,
            I => \Lab_UT.didp.Stens_subtractor.q_RNI775L5_0Z0Z_3\
        );

    \I__6146\ : CascadeMux
    port map (
            O => \N__26605\,
            I => \Lab_UT.didp.Stens_subtractor.q_RNI775L5_0Z0Z_3_cascade_\
        );

    \I__6145\ : CascadeMux
    port map (
            O => \N__26602\,
            I => \N__26599\
        );

    \I__6144\ : InMux
    port map (
            O => \N__26599\,
            I => \N__26596\
        );

    \I__6143\ : LocalMux
    port map (
            O => \N__26596\,
            I => \N__26593\
        );

    \I__6142\ : Odrv4
    port map (
            O => \N__26593\,
            I => \Lab_UT.didp.Stens_subtractor.un1_q_c2\
        );

    \I__6141\ : InMux
    port map (
            O => \N__26590\,
            I => \N__26587\
        );

    \I__6140\ : LocalMux
    port map (
            O => \N__26587\,
            I => \N__26584\
        );

    \I__6139\ : Span4Mux_v
    port map (
            O => \N__26584\,
            I => \N__26580\
        );

    \I__6138\ : InMux
    port map (
            O => \N__26583\,
            I => \N__26577\
        );

    \I__6137\ : IoSpan4Mux
    port map (
            O => \N__26580\,
            I => \N__26572\
        );

    \I__6136\ : LocalMux
    port map (
            O => \N__26577\,
            I => \N__26572\
        );

    \I__6135\ : Odrv4
    port map (
            O => \N__26572\,
            I => \Lab_UT.didp.Stens_subtractor.q_RNI8PD76Z0Z_1\
        );

    \I__6134\ : InMux
    port map (
            O => \N__26569\,
            I => \N__26566\
        );

    \I__6133\ : LocalMux
    port map (
            O => \N__26566\,
            I => \N__26562\
        );

    \I__6132\ : InMux
    port map (
            O => \N__26565\,
            I => \N__26559\
        );

    \I__6131\ : Span4Mux_v
    port map (
            O => \N__26562\,
            I => \N__26554\
        );

    \I__6130\ : LocalMux
    port map (
            O => \N__26559\,
            I => \N__26554\
        );

    \I__6129\ : Odrv4
    port map (
            O => \N__26554\,
            I => \Lab_UT.ld_enable_Stens\
        );

    \I__6128\ : InMux
    port map (
            O => \N__26551\,
            I => \N__26548\
        );

    \I__6127\ : LocalMux
    port map (
            O => \N__26548\,
            I => \N__26545\
        );

    \I__6126\ : Odrv4
    port map (
            O => \N__26545\,
            I => \Lab_UT.didp.Stens_subtractor.q_7_i_1_1\
        );

    \I__6125\ : InMux
    port map (
            O => \N__26542\,
            I => \N__26537\
        );

    \I__6124\ : InMux
    port map (
            O => \N__26541\,
            I => \N__26532\
        );

    \I__6123\ : InMux
    port map (
            O => \N__26540\,
            I => \N__26532\
        );

    \I__6122\ : LocalMux
    port map (
            O => \N__26537\,
            I => \N__26527\
        );

    \I__6121\ : LocalMux
    port map (
            O => \N__26532\,
            I => \N__26527\
        );

    \I__6120\ : Span4Mux_h
    port map (
            O => \N__26527\,
            I => \N__26523\
        );

    \I__6119\ : InMux
    port map (
            O => \N__26526\,
            I => \N__26520\
        );

    \I__6118\ : Odrv4
    port map (
            O => \N__26523\,
            I => \Lab_UT.display.N_152\
        );

    \I__6117\ : LocalMux
    port map (
            O => \N__26520\,
            I => \Lab_UT.display.N_152\
        );

    \I__6116\ : CascadeMux
    port map (
            O => \N__26515\,
            I => \N__26512\
        );

    \I__6115\ : InMux
    port map (
            O => \N__26512\,
            I => \N__26504\
        );

    \I__6114\ : InMux
    port map (
            O => \N__26511\,
            I => \N__26504\
        );

    \I__6113\ : CascadeMux
    port map (
            O => \N__26510\,
            I => \N__26497\
        );

    \I__6112\ : InMux
    port map (
            O => \N__26509\,
            I => \N__26492\
        );

    \I__6111\ : LocalMux
    port map (
            O => \N__26504\,
            I => \N__26487\
        );

    \I__6110\ : InMux
    port map (
            O => \N__26503\,
            I => \N__26483\
        );

    \I__6109\ : InMux
    port map (
            O => \N__26502\,
            I => \N__26478\
        );

    \I__6108\ : InMux
    port map (
            O => \N__26501\,
            I => \N__26478\
        );

    \I__6107\ : InMux
    port map (
            O => \N__26500\,
            I => \N__26469\
        );

    \I__6106\ : InMux
    port map (
            O => \N__26497\,
            I => \N__26469\
        );

    \I__6105\ : InMux
    port map (
            O => \N__26496\,
            I => \N__26469\
        );

    \I__6104\ : InMux
    port map (
            O => \N__26495\,
            I => \N__26469\
        );

    \I__6103\ : LocalMux
    port map (
            O => \N__26492\,
            I => \N__26466\
        );

    \I__6102\ : InMux
    port map (
            O => \N__26491\,
            I => \N__26461\
        );

    \I__6101\ : InMux
    port map (
            O => \N__26490\,
            I => \N__26461\
        );

    \I__6100\ : Span4Mux_h
    port map (
            O => \N__26487\,
            I => \N__26458\
        );

    \I__6099\ : InMux
    port map (
            O => \N__26486\,
            I => \N__26455\
        );

    \I__6098\ : LocalMux
    port map (
            O => \N__26483\,
            I => \Lab_UT.display.cntZ0Z_1\
        );

    \I__6097\ : LocalMux
    port map (
            O => \N__26478\,
            I => \Lab_UT.display.cntZ0Z_1\
        );

    \I__6096\ : LocalMux
    port map (
            O => \N__26469\,
            I => \Lab_UT.display.cntZ0Z_1\
        );

    \I__6095\ : Odrv4
    port map (
            O => \N__26466\,
            I => \Lab_UT.display.cntZ0Z_1\
        );

    \I__6094\ : LocalMux
    port map (
            O => \N__26461\,
            I => \Lab_UT.display.cntZ0Z_1\
        );

    \I__6093\ : Odrv4
    port map (
            O => \N__26458\,
            I => \Lab_UT.display.cntZ0Z_1\
        );

    \I__6092\ : LocalMux
    port map (
            O => \N__26455\,
            I => \Lab_UT.display.cntZ0Z_1\
        );

    \I__6091\ : InMux
    port map (
            O => \N__26440\,
            I => \N__26434\
        );

    \I__6090\ : InMux
    port map (
            O => \N__26439\,
            I => \N__26434\
        );

    \I__6089\ : LocalMux
    port map (
            O => \N__26434\,
            I => \N__26431\
        );

    \I__6088\ : Odrv4
    port map (
            O => \N__26431\,
            I => \Lab_UT.display.N_92\
        );

    \I__6087\ : InMux
    port map (
            O => \N__26428\,
            I => \N__26418\
        );

    \I__6086\ : InMux
    port map (
            O => \N__26427\,
            I => \N__26418\
        );

    \I__6085\ : InMux
    port map (
            O => \N__26426\,
            I => \N__26418\
        );

    \I__6084\ : InMux
    port map (
            O => \N__26425\,
            I => \N__26414\
        );

    \I__6083\ : LocalMux
    port map (
            O => \N__26418\,
            I => \N__26411\
        );

    \I__6082\ : CascadeMux
    port map (
            O => \N__26417\,
            I => \N__26403\
        );

    \I__6081\ : LocalMux
    port map (
            O => \N__26414\,
            I => \N__26398\
        );

    \I__6080\ : Span4Mux_h
    port map (
            O => \N__26411\,
            I => \N__26395\
        );

    \I__6079\ : InMux
    port map (
            O => \N__26410\,
            I => \N__26386\
        );

    \I__6078\ : InMux
    port map (
            O => \N__26409\,
            I => \N__26386\
        );

    \I__6077\ : InMux
    port map (
            O => \N__26408\,
            I => \N__26386\
        );

    \I__6076\ : InMux
    port map (
            O => \N__26407\,
            I => \N__26386\
        );

    \I__6075\ : InMux
    port map (
            O => \N__26406\,
            I => \N__26383\
        );

    \I__6074\ : InMux
    port map (
            O => \N__26403\,
            I => \N__26376\
        );

    \I__6073\ : InMux
    port map (
            O => \N__26402\,
            I => \N__26376\
        );

    \I__6072\ : InMux
    port map (
            O => \N__26401\,
            I => \N__26376\
        );

    \I__6071\ : Odrv4
    port map (
            O => \N__26398\,
            I => \Lab_UT.display.cntZ0Z_2\
        );

    \I__6070\ : Odrv4
    port map (
            O => \N__26395\,
            I => \Lab_UT.display.cntZ0Z_2\
        );

    \I__6069\ : LocalMux
    port map (
            O => \N__26386\,
            I => \Lab_UT.display.cntZ0Z_2\
        );

    \I__6068\ : LocalMux
    port map (
            O => \N__26383\,
            I => \Lab_UT.display.cntZ0Z_2\
        );

    \I__6067\ : LocalMux
    port map (
            O => \N__26376\,
            I => \Lab_UT.display.cntZ0Z_2\
        );

    \I__6066\ : CascadeMux
    port map (
            O => \N__26365\,
            I => \N__26362\
        );

    \I__6065\ : InMux
    port map (
            O => \N__26362\,
            I => \N__26359\
        );

    \I__6064\ : LocalMux
    port map (
            O => \N__26359\,
            I => \N__26356\
        );

    \I__6063\ : Span4Mux_v
    port map (
            O => \N__26356\,
            I => \N__26351\
        );

    \I__6062\ : InMux
    port map (
            O => \N__26355\,
            I => \N__26346\
        );

    \I__6061\ : InMux
    port map (
            O => \N__26354\,
            I => \N__26346\
        );

    \I__6060\ : Odrv4
    port map (
            O => \N__26351\,
            I => \Lab_UT.di_AMtens_1\
        );

    \I__6059\ : LocalMux
    port map (
            O => \N__26346\,
            I => \Lab_UT.di_AMtens_1\
        );

    \I__6058\ : CascadeMux
    port map (
            O => \N__26341\,
            I => \N__26338\
        );

    \I__6057\ : InMux
    port map (
            O => \N__26338\,
            I => \N__26328\
        );

    \I__6056\ : InMux
    port map (
            O => \N__26337\,
            I => \N__26321\
        );

    \I__6055\ : InMux
    port map (
            O => \N__26336\,
            I => \N__26321\
        );

    \I__6054\ : InMux
    port map (
            O => \N__26335\,
            I => \N__26321\
        );

    \I__6053\ : CascadeMux
    port map (
            O => \N__26334\,
            I => \N__26318\
        );

    \I__6052\ : InMux
    port map (
            O => \N__26333\,
            I => \N__26310\
        );

    \I__6051\ : InMux
    port map (
            O => \N__26332\,
            I => \N__26310\
        );

    \I__6050\ : InMux
    port map (
            O => \N__26331\,
            I => \N__26310\
        );

    \I__6049\ : LocalMux
    port map (
            O => \N__26328\,
            I => \N__26305\
        );

    \I__6048\ : LocalMux
    port map (
            O => \N__26321\,
            I => \N__26305\
        );

    \I__6047\ : InMux
    port map (
            O => \N__26318\,
            I => \N__26302\
        );

    \I__6046\ : CascadeMux
    port map (
            O => \N__26317\,
            I => \N__26294\
        );

    \I__6045\ : LocalMux
    port map (
            O => \N__26310\,
            I => \N__26289\
        );

    \I__6044\ : Span4Mux_h
    port map (
            O => \N__26305\,
            I => \N__26284\
        );

    \I__6043\ : LocalMux
    port map (
            O => \N__26302\,
            I => \N__26284\
        );

    \I__6042\ : InMux
    port map (
            O => \N__26301\,
            I => \N__26273\
        );

    \I__6041\ : InMux
    port map (
            O => \N__26300\,
            I => \N__26273\
        );

    \I__6040\ : InMux
    port map (
            O => \N__26299\,
            I => \N__26273\
        );

    \I__6039\ : InMux
    port map (
            O => \N__26298\,
            I => \N__26273\
        );

    \I__6038\ : InMux
    port map (
            O => \N__26297\,
            I => \N__26273\
        );

    \I__6037\ : InMux
    port map (
            O => \N__26294\,
            I => \N__26266\
        );

    \I__6036\ : InMux
    port map (
            O => \N__26293\,
            I => \N__26266\
        );

    \I__6035\ : InMux
    port map (
            O => \N__26292\,
            I => \N__26266\
        );

    \I__6034\ : Odrv4
    port map (
            O => \N__26289\,
            I => \Lab_UT.display.cntZ0Z_0\
        );

    \I__6033\ : Odrv4
    port map (
            O => \N__26284\,
            I => \Lab_UT.display.cntZ0Z_0\
        );

    \I__6032\ : LocalMux
    port map (
            O => \N__26273\,
            I => \Lab_UT.display.cntZ0Z_0\
        );

    \I__6031\ : LocalMux
    port map (
            O => \N__26266\,
            I => \Lab_UT.display.cntZ0Z_0\
        );

    \I__6030\ : InMux
    port map (
            O => \N__26257\,
            I => \N__26254\
        );

    \I__6029\ : LocalMux
    port map (
            O => \N__26254\,
            I => \N__26251\
        );

    \I__6028\ : Span4Mux_h
    port map (
            O => \N__26251\,
            I => \N__26248\
        );

    \I__6027\ : Odrv4
    port map (
            O => \N__26248\,
            I => \Lab_UT.display.N_112\
        );

    \I__6026\ : CascadeMux
    port map (
            O => \N__26245\,
            I => \Lab_UT.didp.Sones_subtractor.q_RNO_0Z0Z_3_cascade_\
        );

    \I__6025\ : CascadeMux
    port map (
            O => \N__26242\,
            I => \N__26239\
        );

    \I__6024\ : InMux
    port map (
            O => \N__26239\,
            I => \N__26236\
        );

    \I__6023\ : LocalMux
    port map (
            O => \N__26236\,
            I => \Lab_UT.didp.Sones_subtractor.q_RNO_0_0_2\
        );

    \I__6022\ : InMux
    port map (
            O => \N__26233\,
            I => \N__26230\
        );

    \I__6021\ : LocalMux
    port map (
            O => \N__26230\,
            I => \N__26226\
        );

    \I__6020\ : InMux
    port map (
            O => \N__26229\,
            I => \N__26220\
        );

    \I__6019\ : Span4Mux_v
    port map (
            O => \N__26226\,
            I => \N__26217\
        );

    \I__6018\ : InMux
    port map (
            O => \N__26225\,
            I => \N__26214\
        );

    \I__6017\ : InMux
    port map (
            O => \N__26224\,
            I => \N__26209\
        );

    \I__6016\ : InMux
    port map (
            O => \N__26223\,
            I => \N__26209\
        );

    \I__6015\ : LocalMux
    port map (
            O => \N__26220\,
            I => \N__26206\
        );

    \I__6014\ : Odrv4
    port map (
            O => \N__26217\,
            I => \Lab_UT.didp.di_Sones_2\
        );

    \I__6013\ : LocalMux
    port map (
            O => \N__26214\,
            I => \Lab_UT.didp.di_Sones_2\
        );

    \I__6012\ : LocalMux
    port map (
            O => \N__26209\,
            I => \Lab_UT.didp.di_Sones_2\
        );

    \I__6011\ : Odrv4
    port map (
            O => \N__26206\,
            I => \Lab_UT.didp.di_Sones_2\
        );

    \I__6010\ : InMux
    port map (
            O => \N__26197\,
            I => \N__26194\
        );

    \I__6009\ : LocalMux
    port map (
            O => \N__26194\,
            I => \N__26189\
        );

    \I__6008\ : CascadeMux
    port map (
            O => \N__26193\,
            I => \N__26185\
        );

    \I__6007\ : CascadeMux
    port map (
            O => \N__26192\,
            I => \N__26182\
        );

    \I__6006\ : Span4Mux_v
    port map (
            O => \N__26189\,
            I => \N__26179\
        );

    \I__6005\ : InMux
    port map (
            O => \N__26188\,
            I => \N__26176\
        );

    \I__6004\ : InMux
    port map (
            O => \N__26185\,
            I => \N__26171\
        );

    \I__6003\ : InMux
    port map (
            O => \N__26182\,
            I => \N__26171\
        );

    \I__6002\ : Sp12to4
    port map (
            O => \N__26179\,
            I => \N__26166\
        );

    \I__6001\ : LocalMux
    port map (
            O => \N__26176\,
            I => \N__26166\
        );

    \I__6000\ : LocalMux
    port map (
            O => \N__26171\,
            I => \Lab_UT.didp.di_Sones_3\
        );

    \I__5999\ : Odrv12
    port map (
            O => \N__26166\,
            I => \Lab_UT.didp.di_Sones_3\
        );

    \I__5998\ : CascadeMux
    port map (
            O => \N__26161\,
            I => \Lab_UT.didp.Sones_subtractor.un8_Mtens_ce_cascade_\
        );

    \I__5997\ : CascadeMux
    port map (
            O => \N__26158\,
            I => \N__26153\
        );

    \I__5996\ : InMux
    port map (
            O => \N__26157\,
            I => \N__26138\
        );

    \I__5995\ : InMux
    port map (
            O => \N__26156\,
            I => \N__26138\
        );

    \I__5994\ : InMux
    port map (
            O => \N__26153\,
            I => \N__26135\
        );

    \I__5993\ : InMux
    port map (
            O => \N__26152\,
            I => \N__26130\
        );

    \I__5992\ : InMux
    port map (
            O => \N__26151\,
            I => \N__26130\
        );

    \I__5991\ : InMux
    port map (
            O => \N__26150\,
            I => \N__26127\
        );

    \I__5990\ : InMux
    port map (
            O => \N__26149\,
            I => \N__26124\
        );

    \I__5989\ : InMux
    port map (
            O => \N__26148\,
            I => \N__26121\
        );

    \I__5988\ : InMux
    port map (
            O => \N__26147\,
            I => \N__26118\
        );

    \I__5987\ : InMux
    port map (
            O => \N__26146\,
            I => \N__26115\
        );

    \I__5986\ : InMux
    port map (
            O => \N__26145\,
            I => \N__26110\
        );

    \I__5985\ : InMux
    port map (
            O => \N__26144\,
            I => \N__26110\
        );

    \I__5984\ : InMux
    port map (
            O => \N__26143\,
            I => \N__26107\
        );

    \I__5983\ : LocalMux
    port map (
            O => \N__26138\,
            I => \N__26060\
        );

    \I__5982\ : LocalMux
    port map (
            O => \N__26135\,
            I => \N__26057\
        );

    \I__5981\ : LocalMux
    port map (
            O => \N__26130\,
            I => \N__26054\
        );

    \I__5980\ : LocalMux
    port map (
            O => \N__26127\,
            I => \N__26051\
        );

    \I__5979\ : LocalMux
    port map (
            O => \N__26124\,
            I => \N__26034\
        );

    \I__5978\ : LocalMux
    port map (
            O => \N__26121\,
            I => \N__26031\
        );

    \I__5977\ : LocalMux
    port map (
            O => \N__26118\,
            I => \N__26028\
        );

    \I__5976\ : LocalMux
    port map (
            O => \N__26115\,
            I => \N__26025\
        );

    \I__5975\ : LocalMux
    port map (
            O => \N__26110\,
            I => \N__26022\
        );

    \I__5974\ : LocalMux
    port map (
            O => \N__26107\,
            I => \N__26019\
        );

    \I__5973\ : SRMux
    port map (
            O => \N__26106\,
            I => \N__25882\
        );

    \I__5972\ : SRMux
    port map (
            O => \N__26105\,
            I => \N__25882\
        );

    \I__5971\ : SRMux
    port map (
            O => \N__26104\,
            I => \N__25882\
        );

    \I__5970\ : SRMux
    port map (
            O => \N__26103\,
            I => \N__25882\
        );

    \I__5969\ : SRMux
    port map (
            O => \N__26102\,
            I => \N__25882\
        );

    \I__5968\ : SRMux
    port map (
            O => \N__26101\,
            I => \N__25882\
        );

    \I__5967\ : SRMux
    port map (
            O => \N__26100\,
            I => \N__25882\
        );

    \I__5966\ : SRMux
    port map (
            O => \N__26099\,
            I => \N__25882\
        );

    \I__5965\ : SRMux
    port map (
            O => \N__26098\,
            I => \N__25882\
        );

    \I__5964\ : SRMux
    port map (
            O => \N__26097\,
            I => \N__25882\
        );

    \I__5963\ : SRMux
    port map (
            O => \N__26096\,
            I => \N__25882\
        );

    \I__5962\ : SRMux
    port map (
            O => \N__26095\,
            I => \N__25882\
        );

    \I__5961\ : SRMux
    port map (
            O => \N__26094\,
            I => \N__25882\
        );

    \I__5960\ : SRMux
    port map (
            O => \N__26093\,
            I => \N__25882\
        );

    \I__5959\ : SRMux
    port map (
            O => \N__26092\,
            I => \N__25882\
        );

    \I__5958\ : SRMux
    port map (
            O => \N__26091\,
            I => \N__25882\
        );

    \I__5957\ : SRMux
    port map (
            O => \N__26090\,
            I => \N__25882\
        );

    \I__5956\ : SRMux
    port map (
            O => \N__26089\,
            I => \N__25882\
        );

    \I__5955\ : SRMux
    port map (
            O => \N__26088\,
            I => \N__25882\
        );

    \I__5954\ : SRMux
    port map (
            O => \N__26087\,
            I => \N__25882\
        );

    \I__5953\ : SRMux
    port map (
            O => \N__26086\,
            I => \N__25882\
        );

    \I__5952\ : SRMux
    port map (
            O => \N__26085\,
            I => \N__25882\
        );

    \I__5951\ : SRMux
    port map (
            O => \N__26084\,
            I => \N__25882\
        );

    \I__5950\ : SRMux
    port map (
            O => \N__26083\,
            I => \N__25882\
        );

    \I__5949\ : SRMux
    port map (
            O => \N__26082\,
            I => \N__25882\
        );

    \I__5948\ : SRMux
    port map (
            O => \N__26081\,
            I => \N__25882\
        );

    \I__5947\ : SRMux
    port map (
            O => \N__26080\,
            I => \N__25882\
        );

    \I__5946\ : SRMux
    port map (
            O => \N__26079\,
            I => \N__25882\
        );

    \I__5945\ : SRMux
    port map (
            O => \N__26078\,
            I => \N__25882\
        );

    \I__5944\ : SRMux
    port map (
            O => \N__26077\,
            I => \N__25882\
        );

    \I__5943\ : SRMux
    port map (
            O => \N__26076\,
            I => \N__25882\
        );

    \I__5942\ : SRMux
    port map (
            O => \N__26075\,
            I => \N__25882\
        );

    \I__5941\ : SRMux
    port map (
            O => \N__26074\,
            I => \N__25882\
        );

    \I__5940\ : SRMux
    port map (
            O => \N__26073\,
            I => \N__25882\
        );

    \I__5939\ : SRMux
    port map (
            O => \N__26072\,
            I => \N__25882\
        );

    \I__5938\ : SRMux
    port map (
            O => \N__26071\,
            I => \N__25882\
        );

    \I__5937\ : SRMux
    port map (
            O => \N__26070\,
            I => \N__25882\
        );

    \I__5936\ : SRMux
    port map (
            O => \N__26069\,
            I => \N__25882\
        );

    \I__5935\ : SRMux
    port map (
            O => \N__26068\,
            I => \N__25882\
        );

    \I__5934\ : SRMux
    port map (
            O => \N__26067\,
            I => \N__25882\
        );

    \I__5933\ : SRMux
    port map (
            O => \N__26066\,
            I => \N__25882\
        );

    \I__5932\ : SRMux
    port map (
            O => \N__26065\,
            I => \N__25882\
        );

    \I__5931\ : SRMux
    port map (
            O => \N__26064\,
            I => \N__25882\
        );

    \I__5930\ : SRMux
    port map (
            O => \N__26063\,
            I => \N__25882\
        );

    \I__5929\ : Glb2LocalMux
    port map (
            O => \N__26060\,
            I => \N__25882\
        );

    \I__5928\ : Glb2LocalMux
    port map (
            O => \N__26057\,
            I => \N__25882\
        );

    \I__5927\ : Glb2LocalMux
    port map (
            O => \N__26054\,
            I => \N__25882\
        );

    \I__5926\ : Glb2LocalMux
    port map (
            O => \N__26051\,
            I => \N__25882\
        );

    \I__5925\ : SRMux
    port map (
            O => \N__26050\,
            I => \N__25882\
        );

    \I__5924\ : SRMux
    port map (
            O => \N__26049\,
            I => \N__25882\
        );

    \I__5923\ : SRMux
    port map (
            O => \N__26048\,
            I => \N__25882\
        );

    \I__5922\ : SRMux
    port map (
            O => \N__26047\,
            I => \N__25882\
        );

    \I__5921\ : SRMux
    port map (
            O => \N__26046\,
            I => \N__25882\
        );

    \I__5920\ : SRMux
    port map (
            O => \N__26045\,
            I => \N__25882\
        );

    \I__5919\ : SRMux
    port map (
            O => \N__26044\,
            I => \N__25882\
        );

    \I__5918\ : SRMux
    port map (
            O => \N__26043\,
            I => \N__25882\
        );

    \I__5917\ : SRMux
    port map (
            O => \N__26042\,
            I => \N__25882\
        );

    \I__5916\ : SRMux
    port map (
            O => \N__26041\,
            I => \N__25882\
        );

    \I__5915\ : SRMux
    port map (
            O => \N__26040\,
            I => \N__25882\
        );

    \I__5914\ : SRMux
    port map (
            O => \N__26039\,
            I => \N__25882\
        );

    \I__5913\ : SRMux
    port map (
            O => \N__26038\,
            I => \N__25882\
        );

    \I__5912\ : SRMux
    port map (
            O => \N__26037\,
            I => \N__25882\
        );

    \I__5911\ : Glb2LocalMux
    port map (
            O => \N__26034\,
            I => \N__25882\
        );

    \I__5910\ : Glb2LocalMux
    port map (
            O => \N__26031\,
            I => \N__25882\
        );

    \I__5909\ : Glb2LocalMux
    port map (
            O => \N__26028\,
            I => \N__25882\
        );

    \I__5908\ : Glb2LocalMux
    port map (
            O => \N__26025\,
            I => \N__25882\
        );

    \I__5907\ : Glb2LocalMux
    port map (
            O => \N__26022\,
            I => \N__25882\
        );

    \I__5906\ : Glb2LocalMux
    port map (
            O => \N__26019\,
            I => \N__25882\
        );

    \I__5905\ : GlobalMux
    port map (
            O => \N__25882\,
            I => \N__25879\
        );

    \I__5904\ : gio2CtrlBuf
    port map (
            O => \N__25879\,
            I => rst_g
        );

    \I__5903\ : InMux
    port map (
            O => \N__25876\,
            I => \N__25870\
        );

    \I__5902\ : InMux
    port map (
            O => \N__25875\,
            I => \N__25870\
        );

    \I__5901\ : LocalMux
    port map (
            O => \N__25870\,
            I => \Lab_UT.display.N_106\
        );

    \I__5900\ : InMux
    port map (
            O => \N__25867\,
            I => \N__25862\
        );

    \I__5899\ : InMux
    port map (
            O => \N__25866\,
            I => \N__25857\
        );

    \I__5898\ : InMux
    port map (
            O => \N__25865\,
            I => \N__25857\
        );

    \I__5897\ : LocalMux
    port map (
            O => \N__25862\,
            I => \Lab_UT.display.N_151\
        );

    \I__5896\ : LocalMux
    port map (
            O => \N__25857\,
            I => \Lab_UT.display.N_151\
        );

    \I__5895\ : InMux
    port map (
            O => \N__25852\,
            I => \N__25848\
        );

    \I__5894\ : InMux
    port map (
            O => \N__25851\,
            I => \N__25845\
        );

    \I__5893\ : LocalMux
    port map (
            O => \N__25848\,
            I => \N__25840\
        );

    \I__5892\ : LocalMux
    port map (
            O => \N__25845\,
            I => \N__25837\
        );

    \I__5891\ : InMux
    port map (
            O => \N__25844\,
            I => \N__25834\
        );

    \I__5890\ : InMux
    port map (
            O => \N__25843\,
            I => \N__25831\
        );

    \I__5889\ : Span4Mux_h
    port map (
            O => \N__25840\,
            I => \N__25828\
        );

    \I__5888\ : Span4Mux_s3_h
    port map (
            O => \N__25837\,
            I => \N__25823\
        );

    \I__5887\ : LocalMux
    port map (
            O => \N__25834\,
            I => \N__25823\
        );

    \I__5886\ : LocalMux
    port map (
            O => \N__25831\,
            I => \Lab_UT.di_AMtens_2\
        );

    \I__5885\ : Odrv4
    port map (
            O => \N__25828\,
            I => \Lab_UT.di_AMtens_2\
        );

    \I__5884\ : Odrv4
    port map (
            O => \N__25823\,
            I => \Lab_UT.di_AMtens_2\
        );

    \I__5883\ : InMux
    port map (
            O => \N__25816\,
            I => \N__25813\
        );

    \I__5882\ : LocalMux
    port map (
            O => \N__25813\,
            I => \Lab_UT.display.N_115\
        );

    \I__5881\ : InMux
    port map (
            O => \N__25810\,
            I => \N__25806\
        );

    \I__5880\ : CascadeMux
    port map (
            O => \N__25809\,
            I => \N__25803\
        );

    \I__5879\ : LocalMux
    port map (
            O => \N__25806\,
            I => \N__25799\
        );

    \I__5878\ : InMux
    port map (
            O => \N__25803\,
            I => \N__25796\
        );

    \I__5877\ : InMux
    port map (
            O => \N__25802\,
            I => \N__25793\
        );

    \I__5876\ : Span4Mux_s3_h
    port map (
            O => \N__25799\,
            I => \N__25788\
        );

    \I__5875\ : LocalMux
    port map (
            O => \N__25796\,
            I => \N__25788\
        );

    \I__5874\ : LocalMux
    port map (
            O => \N__25793\,
            I => \Lab_UT.di_AStens_1\
        );

    \I__5873\ : Odrv4
    port map (
            O => \N__25788\,
            I => \Lab_UT.di_AStens_1\
        );

    \I__5872\ : CascadeMux
    port map (
            O => \N__25783\,
            I => \Lab_UT.display.N_108_cascade_\
        );

    \I__5871\ : InMux
    port map (
            O => \N__25780\,
            I => \N__25776\
        );

    \I__5870\ : InMux
    port map (
            O => \N__25779\,
            I => \N__25772\
        );

    \I__5869\ : LocalMux
    port map (
            O => \N__25776\,
            I => \N__25769\
        );

    \I__5868\ : InMux
    port map (
            O => \N__25775\,
            I => \N__25766\
        );

    \I__5867\ : LocalMux
    port map (
            O => \N__25772\,
            I => \N__25763\
        );

    \I__5866\ : Span4Mux_v
    port map (
            O => \N__25769\,
            I => \N__25760\
        );

    \I__5865\ : LocalMux
    port map (
            O => \N__25766\,
            I => \Lab_UT.di_AMones_1\
        );

    \I__5864\ : Odrv4
    port map (
            O => \N__25763\,
            I => \Lab_UT.di_AMones_1\
        );

    \I__5863\ : Odrv4
    port map (
            O => \N__25760\,
            I => \Lab_UT.di_AMones_1\
        );

    \I__5862\ : InMux
    port map (
            O => \N__25753\,
            I => \N__25750\
        );

    \I__5861\ : LocalMux
    port map (
            O => \N__25750\,
            I => \N__25747\
        );

    \I__5860\ : Span4Mux_h
    port map (
            O => \N__25747\,
            I => \N__25744\
        );

    \I__5859\ : Odrv4
    port map (
            O => \N__25744\,
            I => \Lab_UT.display.dOutP_0_iv_i_0_1\
        );

    \I__5858\ : CascadeMux
    port map (
            O => \N__25741\,
            I => \N__25738\
        );

    \I__5857\ : InMux
    port map (
            O => \N__25738\,
            I => \N__25735\
        );

    \I__5856\ : LocalMux
    port map (
            O => \N__25735\,
            I => \Lab_UT.displayAlarmZ0Z_0\
        );

    \I__5855\ : InMux
    port map (
            O => \N__25732\,
            I => \N__25729\
        );

    \I__5854\ : LocalMux
    port map (
            O => \N__25729\,
            I => \N__25725\
        );

    \I__5853\ : InMux
    port map (
            O => \N__25728\,
            I => \N__25721\
        );

    \I__5852\ : Span4Mux_v
    port map (
            O => \N__25725\,
            I => \N__25718\
        );

    \I__5851\ : InMux
    port map (
            O => \N__25724\,
            I => \N__25715\
        );

    \I__5850\ : LocalMux
    port map (
            O => \N__25721\,
            I => \Lab_UT.di_AStens_0\
        );

    \I__5849\ : Odrv4
    port map (
            O => \N__25718\,
            I => \Lab_UT.di_AStens_0\
        );

    \I__5848\ : LocalMux
    port map (
            O => \N__25715\,
            I => \Lab_UT.di_AStens_0\
        );

    \I__5847\ : InMux
    port map (
            O => \N__25708\,
            I => \N__25705\
        );

    \I__5846\ : LocalMux
    port map (
            O => \N__25705\,
            I => \Lab_UT.display.N_130\
        );

    \I__5845\ : CascadeMux
    port map (
            O => \N__25702\,
            I => \Lab_UT.display.dOutP_0_iv_i_0_0_cascade_\
        );

    \I__5844\ : InMux
    port map (
            O => \N__25699\,
            I => \N__25696\
        );

    \I__5843\ : LocalMux
    port map (
            O => \N__25696\,
            I => \N__25693\
        );

    \I__5842\ : Span4Mux_v
    port map (
            O => \N__25693\,
            I => \N__25690\
        );

    \I__5841\ : Odrv4
    port map (
            O => \N__25690\,
            I => \Lab_UT.display.dOutP_0_iv_i_1_0\
        );

    \I__5840\ : CascadeMux
    port map (
            O => \N__25687\,
            I => \N__25684\
        );

    \I__5839\ : InMux
    port map (
            O => \N__25684\,
            I => \N__25677\
        );

    \I__5838\ : InMux
    port map (
            O => \N__25683\,
            I => \N__25677\
        );

    \I__5837\ : InMux
    port map (
            O => \N__25682\,
            I => \N__25674\
        );

    \I__5836\ : LocalMux
    port map (
            O => \N__25677\,
            I => \N__25671\
        );

    \I__5835\ : LocalMux
    port map (
            O => \N__25674\,
            I => \N__25668\
        );

    \I__5834\ : Span4Mux_h
    port map (
            O => \N__25671\,
            I => \N__25665\
        );

    \I__5833\ : Odrv12
    port map (
            O => \N__25668\,
            I => \L3_tx_data_0\
        );

    \I__5832\ : Odrv4
    port map (
            O => \N__25665\,
            I => \L3_tx_data_0\
        );

    \I__5831\ : InMux
    port map (
            O => \N__25660\,
            I => \N__25654\
        );

    \I__5830\ : InMux
    port map (
            O => \N__25659\,
            I => \N__25654\
        );

    \I__5829\ : LocalMux
    port map (
            O => \N__25654\,
            I => \N__25651\
        );

    \I__5828\ : Span4Mux_s2_h
    port map (
            O => \N__25651\,
            I => \N__25648\
        );

    \I__5827\ : Odrv4
    port map (
            O => \N__25648\,
            I => \Lab_UT.display.N_153\
        );

    \I__5826\ : CascadeMux
    port map (
            O => \N__25645\,
            I => \N__25642\
        );

    \I__5825\ : InMux
    port map (
            O => \N__25642\,
            I => \N__25639\
        );

    \I__5824\ : LocalMux
    port map (
            O => \N__25639\,
            I => \N__25636\
        );

    \I__5823\ : Odrv4
    port map (
            O => \N__25636\,
            I => \Lab_UT.displayAlarmZ1Z_2\
        );

    \I__5822\ : InMux
    port map (
            O => \N__25633\,
            I => \N__25630\
        );

    \I__5821\ : LocalMux
    port map (
            O => \N__25630\,
            I => \N__25626\
        );

    \I__5820\ : InMux
    port map (
            O => \N__25629\,
            I => \N__25622\
        );

    \I__5819\ : Span4Mux_s2_h
    port map (
            O => \N__25626\,
            I => \N__25619\
        );

    \I__5818\ : InMux
    port map (
            O => \N__25625\,
            I => \N__25616\
        );

    \I__5817\ : LocalMux
    port map (
            O => \N__25622\,
            I => \Lab_UT.di_AStens_2\
        );

    \I__5816\ : Odrv4
    port map (
            O => \N__25619\,
            I => \Lab_UT.di_AStens_2\
        );

    \I__5815\ : LocalMux
    port map (
            O => \N__25616\,
            I => \Lab_UT.di_AStens_2\
        );

    \I__5814\ : CascadeMux
    port map (
            O => \N__25609\,
            I => \Lab_UT.display.dOutP_0_iv_i_0_2_cascade_\
        );

    \I__5813\ : InMux
    port map (
            O => \N__25606\,
            I => \N__25603\
        );

    \I__5812\ : LocalMux
    port map (
            O => \N__25603\,
            I => \N__25600\
        );

    \I__5811\ : Span4Mux_v
    port map (
            O => \N__25600\,
            I => \N__25597\
        );

    \I__5810\ : Odrv4
    port map (
            O => \N__25597\,
            I => \Lab_UT.display.dOutP_0_iv_i_1_2\
        );

    \I__5809\ : CascadeMux
    port map (
            O => \N__25594\,
            I => \N__25591\
        );

    \I__5808\ : InMux
    port map (
            O => \N__25591\,
            I => \N__25587\
        );

    \I__5807\ : InMux
    port map (
            O => \N__25590\,
            I => \N__25583\
        );

    \I__5806\ : LocalMux
    port map (
            O => \N__25587\,
            I => \N__25580\
        );

    \I__5805\ : InMux
    port map (
            O => \N__25586\,
            I => \N__25577\
        );

    \I__5804\ : LocalMux
    port map (
            O => \N__25583\,
            I => \N__25570\
        );

    \I__5803\ : Span4Mux_s3_v
    port map (
            O => \N__25580\,
            I => \N__25570\
        );

    \I__5802\ : LocalMux
    port map (
            O => \N__25577\,
            I => \N__25570\
        );

    \I__5801\ : Odrv4
    port map (
            O => \N__25570\,
            I => \L3_tx_data_2\
        );

    \I__5800\ : InMux
    port map (
            O => \N__25567\,
            I => \N__25558\
        );

    \I__5799\ : InMux
    port map (
            O => \N__25566\,
            I => \N__25558\
        );

    \I__5798\ : InMux
    port map (
            O => \N__25565\,
            I => \N__25558\
        );

    \I__5797\ : LocalMux
    port map (
            O => \N__25558\,
            I => \N__25555\
        );

    \I__5796\ : Odrv4
    port map (
            O => \N__25555\,
            I => \Lab_UT.display.un42_dOutP_1\
        );

    \I__5795\ : InMux
    port map (
            O => \N__25552\,
            I => \N__25546\
        );

    \I__5794\ : InMux
    port map (
            O => \N__25551\,
            I => \N__25546\
        );

    \I__5793\ : LocalMux
    port map (
            O => \N__25546\,
            I => \N__25543\
        );

    \I__5792\ : Span4Mux_v
    port map (
            O => \N__25543\,
            I => \N__25540\
        );

    \I__5791\ : Odrv4
    port map (
            O => \N__25540\,
            I => \Lab_UT.display.cnt_RNI1STE1Z0Z_1\
        );

    \I__5790\ : CascadeMux
    port map (
            O => \N__25537\,
            I => \Lab_UT.display.N_151_cascade_\
        );

    \I__5789\ : InMux
    port map (
            O => \N__25534\,
            I => \N__25530\
        );

    \I__5788\ : InMux
    port map (
            O => \N__25533\,
            I => \N__25527\
        );

    \I__5787\ : LocalMux
    port map (
            O => \N__25530\,
            I => \N__25523\
        );

    \I__5786\ : LocalMux
    port map (
            O => \N__25527\,
            I => \N__25520\
        );

    \I__5785\ : InMux
    port map (
            O => \N__25526\,
            I => \N__25517\
        );

    \I__5784\ : Span4Mux_s2_h
    port map (
            O => \N__25523\,
            I => \N__25514\
        );

    \I__5783\ : Span4Mux_h
    port map (
            O => \N__25520\,
            I => \N__25511\
        );

    \I__5782\ : LocalMux
    port map (
            O => \N__25517\,
            I => \Lab_UT.di_AMtens_3\
        );

    \I__5781\ : Odrv4
    port map (
            O => \N__25514\,
            I => \Lab_UT.di_AMtens_3\
        );

    \I__5780\ : Odrv4
    port map (
            O => \N__25511\,
            I => \Lab_UT.di_AMtens_3\
        );

    \I__5779\ : InMux
    port map (
            O => \N__25504\,
            I => \N__25501\
        );

    \I__5778\ : LocalMux
    port map (
            O => \N__25501\,
            I => \N__25498\
        );

    \I__5777\ : Odrv4
    port map (
            O => \N__25498\,
            I => \Lab_UT.display.N_124\
        );

    \I__5776\ : CascadeMux
    port map (
            O => \N__25495\,
            I => \Lab_UT.dictrl.decoder.de_littleNZ0Z_1_cascade_\
        );

    \I__5775\ : InMux
    port map (
            O => \N__25492\,
            I => \N__25486\
        );

    \I__5774\ : InMux
    port map (
            O => \N__25491\,
            I => \N__25479\
        );

    \I__5773\ : InMux
    port map (
            O => \N__25490\,
            I => \N__25479\
        );

    \I__5772\ : InMux
    port map (
            O => \N__25489\,
            I => \N__25479\
        );

    \I__5771\ : LocalMux
    port map (
            O => \N__25486\,
            I => \N__25474\
        );

    \I__5770\ : LocalMux
    port map (
            O => \N__25479\,
            I => \N__25471\
        );

    \I__5769\ : InMux
    port map (
            O => \N__25478\,
            I => \N__25466\
        );

    \I__5768\ : InMux
    port map (
            O => \N__25477\,
            I => \N__25466\
        );

    \I__5767\ : Span4Mux_v
    port map (
            O => \N__25474\,
            I => \N__25461\
        );

    \I__5766\ : Span4Mux_v
    port map (
            O => \N__25471\,
            I => \N__25461\
        );

    \I__5765\ : LocalMux
    port map (
            O => \N__25466\,
            I => \Lab_UT_dictrl_decoder_de_cr_2\
        );

    \I__5764\ : Odrv4
    port map (
            O => \N__25461\,
            I => \Lab_UT_dictrl_decoder_de_cr_2\
        );

    \I__5763\ : CascadeMux
    port map (
            O => \N__25456\,
            I => \N__25453\
        );

    \I__5762\ : InMux
    port map (
            O => \N__25453\,
            I => \N__25447\
        );

    \I__5761\ : InMux
    port map (
            O => \N__25452\,
            I => \N__25447\
        );

    \I__5760\ : LocalMux
    port map (
            O => \N__25447\,
            I => \N__25444\
        );

    \I__5759\ : Span4Mux_v
    port map (
            O => \N__25444\,
            I => \N__25441\
        );

    \I__5758\ : Span4Mux_v
    port map (
            O => \N__25441\,
            I => \N__25438\
        );

    \I__5757\ : Odrv4
    port map (
            O => \N__25438\,
            I => \Lab_UT.n_rdy\
        );

    \I__5756\ : InMux
    port map (
            O => \N__25435\,
            I => \N__25432\
        );

    \I__5755\ : LocalMux
    port map (
            O => \N__25432\,
            I => \resetGen.escKeyZ0Z_3\
        );

    \I__5754\ : CEMux
    port map (
            O => \N__25429\,
            I => \N__25408\
        );

    \I__5753\ : CEMux
    port map (
            O => \N__25428\,
            I => \N__25408\
        );

    \I__5752\ : CEMux
    port map (
            O => \N__25427\,
            I => \N__25408\
        );

    \I__5751\ : CEMux
    port map (
            O => \N__25426\,
            I => \N__25408\
        );

    \I__5750\ : CEMux
    port map (
            O => \N__25425\,
            I => \N__25408\
        );

    \I__5749\ : CEMux
    port map (
            O => \N__25424\,
            I => \N__25408\
        );

    \I__5748\ : CEMux
    port map (
            O => \N__25423\,
            I => \N__25408\
        );

    \I__5747\ : GlobalMux
    port map (
            O => \N__25408\,
            I => \N__25405\
        );

    \I__5746\ : gio2CtrlBuf
    port map (
            O => \N__25405\,
            I => \buart.Z_rx.sample_g\
        );

    \I__5745\ : InMux
    port map (
            O => \N__25402\,
            I => \N__25399\
        );

    \I__5744\ : LocalMux
    port map (
            O => \N__25399\,
            I => \N__25391\
        );

    \I__5743\ : InMux
    port map (
            O => \N__25398\,
            I => \N__25386\
        );

    \I__5742\ : InMux
    port map (
            O => \N__25397\,
            I => \N__25386\
        );

    \I__5741\ : InMux
    port map (
            O => \N__25396\,
            I => \N__25381\
        );

    \I__5740\ : InMux
    port map (
            O => \N__25395\,
            I => \N__25381\
        );

    \I__5739\ : InMux
    port map (
            O => \N__25394\,
            I => \N__25378\
        );

    \I__5738\ : Span4Mux_s3_h
    port map (
            O => \N__25391\,
            I => \N__25363\
        );

    \I__5737\ : LocalMux
    port map (
            O => \N__25386\,
            I => \N__25363\
        );

    \I__5736\ : LocalMux
    port map (
            O => \N__25381\,
            I => \N__25363\
        );

    \I__5735\ : LocalMux
    port map (
            O => \N__25378\,
            I => \N__25363\
        );

    \I__5734\ : InMux
    port map (
            O => \N__25377\,
            I => \N__25360\
        );

    \I__5733\ : InMux
    port map (
            O => \N__25376\,
            I => \N__25357\
        );

    \I__5732\ : InMux
    port map (
            O => \N__25375\,
            I => \N__25350\
        );

    \I__5731\ : InMux
    port map (
            O => \N__25374\,
            I => \N__25350\
        );

    \I__5730\ : InMux
    port map (
            O => \N__25373\,
            I => \N__25350\
        );

    \I__5729\ : InMux
    port map (
            O => \N__25372\,
            I => \N__25347\
        );

    \I__5728\ : Span4Mux_h
    port map (
            O => \N__25363\,
            I => \N__25341\
        );

    \I__5727\ : LocalMux
    port map (
            O => \N__25360\,
            I => \N__25334\
        );

    \I__5726\ : LocalMux
    port map (
            O => \N__25357\,
            I => \N__25334\
        );

    \I__5725\ : LocalMux
    port map (
            O => \N__25350\,
            I => \N__25334\
        );

    \I__5724\ : LocalMux
    port map (
            O => \N__25347\,
            I => \N__25331\
        );

    \I__5723\ : InMux
    port map (
            O => \N__25346\,
            I => \N__25324\
        );

    \I__5722\ : InMux
    port map (
            O => \N__25345\,
            I => \N__25324\
        );

    \I__5721\ : InMux
    port map (
            O => \N__25344\,
            I => \N__25324\
        );

    \I__5720\ : Odrv4
    port map (
            O => \N__25341\,
            I => bu_rx_data_7
        );

    \I__5719\ : Odrv12
    port map (
            O => \N__25334\,
            I => bu_rx_data_7
        );

    \I__5718\ : Odrv4
    port map (
            O => \N__25331\,
            I => bu_rx_data_7
        );

    \I__5717\ : LocalMux
    port map (
            O => \N__25324\,
            I => bu_rx_data_7
        );

    \I__5716\ : InMux
    port map (
            O => \N__25315\,
            I => \N__25308\
        );

    \I__5715\ : InMux
    port map (
            O => \N__25314\,
            I => \N__25308\
        );

    \I__5714\ : InMux
    port map (
            O => \N__25313\,
            I => \N__25305\
        );

    \I__5713\ : LocalMux
    port map (
            O => \N__25308\,
            I => \N__25297\
        );

    \I__5712\ : LocalMux
    port map (
            O => \N__25305\,
            I => \N__25294\
        );

    \I__5711\ : InMux
    port map (
            O => \N__25304\,
            I => \N__25291\
        );

    \I__5710\ : InMux
    port map (
            O => \N__25303\,
            I => \N__25288\
        );

    \I__5709\ : InMux
    port map (
            O => \N__25302\,
            I => \N__25283\
        );

    \I__5708\ : InMux
    port map (
            O => \N__25301\,
            I => \N__25283\
        );

    \I__5707\ : InMux
    port map (
            O => \N__25300\,
            I => \N__25280\
        );

    \I__5706\ : Span4Mux_v
    port map (
            O => \N__25297\,
            I => \N__25274\
        );

    \I__5705\ : Span4Mux_s2_v
    port map (
            O => \N__25294\,
            I => \N__25274\
        );

    \I__5704\ : LocalMux
    port map (
            O => \N__25291\,
            I => \N__25269\
        );

    \I__5703\ : LocalMux
    port map (
            O => \N__25288\,
            I => \N__25266\
        );

    \I__5702\ : LocalMux
    port map (
            O => \N__25283\,
            I => \N__25261\
        );

    \I__5701\ : LocalMux
    port map (
            O => \N__25280\,
            I => \N__25261\
        );

    \I__5700\ : InMux
    port map (
            O => \N__25279\,
            I => \N__25257\
        );

    \I__5699\ : Span4Mux_h
    port map (
            O => \N__25274\,
            I => \N__25254\
        );

    \I__5698\ : InMux
    port map (
            O => \N__25273\,
            I => \N__25251\
        );

    \I__5697\ : InMux
    port map (
            O => \N__25272\,
            I => \N__25248\
        );

    \I__5696\ : Span4Mux_v
    port map (
            O => \N__25269\,
            I => \N__25241\
        );

    \I__5695\ : Span4Mux_h
    port map (
            O => \N__25266\,
            I => \N__25241\
        );

    \I__5694\ : Span4Mux_s2_v
    port map (
            O => \N__25261\,
            I => \N__25241\
        );

    \I__5693\ : InMux
    port map (
            O => \N__25260\,
            I => \N__25238\
        );

    \I__5692\ : LocalMux
    port map (
            O => \N__25257\,
            I => bu_rx_data_4
        );

    \I__5691\ : Odrv4
    port map (
            O => \N__25254\,
            I => bu_rx_data_4
        );

    \I__5690\ : LocalMux
    port map (
            O => \N__25251\,
            I => bu_rx_data_4
        );

    \I__5689\ : LocalMux
    port map (
            O => \N__25248\,
            I => bu_rx_data_4
        );

    \I__5688\ : Odrv4
    port map (
            O => \N__25241\,
            I => bu_rx_data_4
        );

    \I__5687\ : LocalMux
    port map (
            O => \N__25238\,
            I => bu_rx_data_4
        );

    \I__5686\ : InMux
    port map (
            O => \N__25225\,
            I => \N__25222\
        );

    \I__5685\ : LocalMux
    port map (
            O => \N__25222\,
            I => \N__25219\
        );

    \I__5684\ : Odrv4
    port map (
            O => \N__25219\,
            I => \Lab_UT.dictrl.decoder.de_atSignZ0Z_5\
        );

    \I__5683\ : CascadeMux
    port map (
            O => \N__25216\,
            I => \N__25213\
        );

    \I__5682\ : InMux
    port map (
            O => \N__25213\,
            I => \N__25201\
        );

    \I__5681\ : InMux
    port map (
            O => \N__25212\,
            I => \N__25201\
        );

    \I__5680\ : InMux
    port map (
            O => \N__25211\,
            I => \N__25201\
        );

    \I__5679\ : InMux
    port map (
            O => \N__25210\,
            I => \N__25201\
        );

    \I__5678\ : LocalMux
    port map (
            O => \N__25201\,
            I => \N__25196\
        );

    \I__5677\ : InMux
    port map (
            O => \N__25200\,
            I => \N__25193\
        );

    \I__5676\ : InMux
    port map (
            O => \N__25199\,
            I => \N__25190\
        );

    \I__5675\ : Sp12to4
    port map (
            O => \N__25196\,
            I => \N__25185\
        );

    \I__5674\ : LocalMux
    port map (
            O => \N__25193\,
            I => \N__25185\
        );

    \I__5673\ : LocalMux
    port map (
            O => \N__25190\,
            I => \Lab_UT.uu0.l_precountZ0Z_0\
        );

    \I__5672\ : Odrv12
    port map (
            O => \N__25185\,
            I => \Lab_UT.uu0.l_precountZ0Z_0\
        );

    \I__5671\ : InMux
    port map (
            O => \N__25180\,
            I => \N__25176\
        );

    \I__5670\ : InMux
    port map (
            O => \N__25179\,
            I => \N__25173\
        );

    \I__5669\ : LocalMux
    port map (
            O => \N__25176\,
            I => \N__25170\
        );

    \I__5668\ : LocalMux
    port map (
            O => \N__25173\,
            I => \N__25167\
        );

    \I__5667\ : Span4Mux_v
    port map (
            O => \N__25170\,
            I => \N__25162\
        );

    \I__5666\ : Span4Mux_s2_h
    port map (
            O => \N__25167\,
            I => \N__25162\
        );

    \I__5665\ : Span4Mux_h
    port map (
            O => \N__25162\,
            I => \N__25157\
        );

    \I__5664\ : InMux
    port map (
            O => \N__25161\,
            I => \N__25152\
        );

    \I__5663\ : InMux
    port map (
            O => \N__25160\,
            I => \N__25152\
        );

    \I__5662\ : Odrv4
    port map (
            O => \N__25157\,
            I => \uu2.un404_ci_0\
        );

    \I__5661\ : LocalMux
    port map (
            O => \N__25152\,
            I => \uu2.un404_ci_0\
        );

    \I__5660\ : InMux
    port map (
            O => \N__25147\,
            I => \N__25143\
        );

    \I__5659\ : InMux
    port map (
            O => \N__25146\,
            I => \N__25140\
        );

    \I__5658\ : LocalMux
    port map (
            O => \N__25143\,
            I => \N__25137\
        );

    \I__5657\ : LocalMux
    port map (
            O => \N__25140\,
            I => \N__25134\
        );

    \I__5656\ : Span4Mux_v
    port map (
            O => \N__25137\,
            I => \N__25126\
        );

    \I__5655\ : Span4Mux_s3_h
    port map (
            O => \N__25134\,
            I => \N__25126\
        );

    \I__5654\ : InMux
    port map (
            O => \N__25133\,
            I => \N__25119\
        );

    \I__5653\ : InMux
    port map (
            O => \N__25132\,
            I => \N__25119\
        );

    \I__5652\ : InMux
    port map (
            O => \N__25131\,
            I => \N__25119\
        );

    \I__5651\ : Odrv4
    port map (
            O => \N__25126\,
            I => \uu2.trig_rd_is_det\
        );

    \I__5650\ : LocalMux
    port map (
            O => \N__25119\,
            I => \uu2.trig_rd_is_det\
        );

    \I__5649\ : CascadeMux
    port map (
            O => \N__25114\,
            I => \N__25111\
        );

    \I__5648\ : InMux
    port map (
            O => \N__25111\,
            I => \N__25105\
        );

    \I__5647\ : InMux
    port map (
            O => \N__25110\,
            I => \N__25100\
        );

    \I__5646\ : InMux
    port map (
            O => \N__25109\,
            I => \N__25100\
        );

    \I__5645\ : InMux
    port map (
            O => \N__25108\,
            I => \N__25097\
        );

    \I__5644\ : LocalMux
    port map (
            O => \N__25105\,
            I => \N__25092\
        );

    \I__5643\ : LocalMux
    port map (
            O => \N__25100\,
            I => \N__25092\
        );

    \I__5642\ : LocalMux
    port map (
            O => \N__25097\,
            I => \N__25089\
        );

    \I__5641\ : Span4Mux_h
    port map (
            O => \N__25092\,
            I => \N__25085\
        );

    \I__5640\ : Span4Mux_h
    port map (
            O => \N__25089\,
            I => \N__25082\
        );

    \I__5639\ : InMux
    port map (
            O => \N__25088\,
            I => \N__25079\
        );

    \I__5638\ : Span4Mux_h
    port map (
            O => \N__25085\,
            I => \N__25076\
        );

    \I__5637\ : Odrv4
    port map (
            O => \N__25082\,
            I => \uu2.r_addrZ0Z_4\
        );

    \I__5636\ : LocalMux
    port map (
            O => \N__25079\,
            I => \uu2.r_addrZ0Z_4\
        );

    \I__5635\ : Odrv4
    port map (
            O => \N__25076\,
            I => \uu2.r_addrZ0Z_4\
        );

    \I__5634\ : InMux
    port map (
            O => \N__25069\,
            I => \N__25066\
        );

    \I__5633\ : LocalMux
    port map (
            O => \N__25066\,
            I => \N__25063\
        );

    \I__5632\ : Span12Mux_s8_v
    port map (
            O => \N__25063\,
            I => \N__25058\
        );

    \I__5631\ : InMux
    port map (
            O => \N__25062\,
            I => \N__25053\
        );

    \I__5630\ : InMux
    port map (
            O => \N__25061\,
            I => \N__25053\
        );

    \I__5629\ : Odrv12
    port map (
            O => \N__25058\,
            I => \Lab_UT.di_AMtens_0\
        );

    \I__5628\ : LocalMux
    port map (
            O => \N__25053\,
            I => \Lab_UT.di_AMtens_0\
        );

    \I__5627\ : CascadeMux
    port map (
            O => \N__25048\,
            I => \N__25042\
        );

    \I__5626\ : CascadeMux
    port map (
            O => \N__25047\,
            I => \N__25036\
        );

    \I__5625\ : CascadeMux
    port map (
            O => \N__25046\,
            I => \N__25033\
        );

    \I__5624\ : InMux
    port map (
            O => \N__25045\,
            I => \N__25026\
        );

    \I__5623\ : InMux
    port map (
            O => \N__25042\,
            I => \N__25026\
        );

    \I__5622\ : InMux
    port map (
            O => \N__25041\,
            I => \N__25026\
        );

    \I__5621\ : InMux
    port map (
            O => \N__25040\,
            I => \N__25016\
        );

    \I__5620\ : CascadeMux
    port map (
            O => \N__25039\,
            I => \N__25013\
        );

    \I__5619\ : InMux
    port map (
            O => \N__25036\,
            I => \N__25005\
        );

    \I__5618\ : InMux
    port map (
            O => \N__25033\,
            I => \N__25002\
        );

    \I__5617\ : LocalMux
    port map (
            O => \N__25026\,
            I => \N__24999\
        );

    \I__5616\ : InMux
    port map (
            O => \N__25025\,
            I => \N__24996\
        );

    \I__5615\ : InMux
    port map (
            O => \N__25024\,
            I => \N__24987\
        );

    \I__5614\ : InMux
    port map (
            O => \N__25023\,
            I => \N__24987\
        );

    \I__5613\ : InMux
    port map (
            O => \N__25022\,
            I => \N__24987\
        );

    \I__5612\ : InMux
    port map (
            O => \N__25021\,
            I => \N__24987\
        );

    \I__5611\ : InMux
    port map (
            O => \N__25020\,
            I => \N__24982\
        );

    \I__5610\ : InMux
    port map (
            O => \N__25019\,
            I => \N__24982\
        );

    \I__5609\ : LocalMux
    port map (
            O => \N__25016\,
            I => \N__24979\
        );

    \I__5608\ : InMux
    port map (
            O => \N__25013\,
            I => \N__24976\
        );

    \I__5607\ : InMux
    port map (
            O => \N__25012\,
            I => \N__24973\
        );

    \I__5606\ : InMux
    port map (
            O => \N__25011\,
            I => \N__24968\
        );

    \I__5605\ : InMux
    port map (
            O => \N__25010\,
            I => \N__24968\
        );

    \I__5604\ : CascadeMux
    port map (
            O => \N__25009\,
            I => \N__24965\
        );

    \I__5603\ : InMux
    port map (
            O => \N__25008\,
            I => \N__24961\
        );

    \I__5602\ : LocalMux
    port map (
            O => \N__25005\,
            I => \N__24958\
        );

    \I__5601\ : LocalMux
    port map (
            O => \N__25002\,
            I => \N__24953\
        );

    \I__5600\ : Span4Mux_s2_h
    port map (
            O => \N__24999\,
            I => \N__24953\
        );

    \I__5599\ : LocalMux
    port map (
            O => \N__24996\,
            I => \N__24950\
        );

    \I__5598\ : LocalMux
    port map (
            O => \N__24987\,
            I => \N__24947\
        );

    \I__5597\ : LocalMux
    port map (
            O => \N__24982\,
            I => \N__24944\
        );

    \I__5596\ : Span4Mux_h
    port map (
            O => \N__24979\,
            I => \N__24935\
        );

    \I__5595\ : LocalMux
    port map (
            O => \N__24976\,
            I => \N__24935\
        );

    \I__5594\ : LocalMux
    port map (
            O => \N__24973\,
            I => \N__24935\
        );

    \I__5593\ : LocalMux
    port map (
            O => \N__24968\,
            I => \N__24935\
        );

    \I__5592\ : InMux
    port map (
            O => \N__24965\,
            I => \N__24930\
        );

    \I__5591\ : InMux
    port map (
            O => \N__24964\,
            I => \N__24930\
        );

    \I__5590\ : LocalMux
    port map (
            O => \N__24961\,
            I => \N__24927\
        );

    \I__5589\ : Span4Mux_h
    port map (
            O => \N__24958\,
            I => \N__24922\
        );

    \I__5588\ : Span4Mux_h
    port map (
            O => \N__24953\,
            I => \N__24922\
        );

    \I__5587\ : Span4Mux_v
    port map (
            O => \N__24950\,
            I => \N__24919\
        );

    \I__5586\ : Span4Mux_v
    port map (
            O => \N__24947\,
            I => \N__24910\
        );

    \I__5585\ : Span4Mux_h
    port map (
            O => \N__24944\,
            I => \N__24910\
        );

    \I__5584\ : Span4Mux_v
    port map (
            O => \N__24935\,
            I => \N__24910\
        );

    \I__5583\ : LocalMux
    port map (
            O => \N__24930\,
            I => \N__24910\
        );

    \I__5582\ : Odrv12
    port map (
            O => \N__24927\,
            I => \Lab_UT.dictrl.currStateZ0Z_2\
        );

    \I__5581\ : Odrv4
    port map (
            O => \N__24922\,
            I => \Lab_UT.dictrl.currStateZ0Z_2\
        );

    \I__5580\ : Odrv4
    port map (
            O => \N__24919\,
            I => \Lab_UT.dictrl.currStateZ0Z_2\
        );

    \I__5579\ : Odrv4
    port map (
            O => \N__24910\,
            I => \Lab_UT.dictrl.currStateZ0Z_2\
        );

    \I__5578\ : CascadeMux
    port map (
            O => \N__24901\,
            I => \N__24894\
        );

    \I__5577\ : CascadeMux
    port map (
            O => \N__24900\,
            I => \N__24891\
        );

    \I__5576\ : CascadeMux
    port map (
            O => \N__24899\,
            I => \N__24882\
        );

    \I__5575\ : CascadeMux
    port map (
            O => \N__24898\,
            I => \N__24879\
        );

    \I__5574\ : CascadeMux
    port map (
            O => \N__24897\,
            I => \N__24875\
        );

    \I__5573\ : InMux
    port map (
            O => \N__24894\,
            I => \N__24871\
        );

    \I__5572\ : InMux
    port map (
            O => \N__24891\,
            I => \N__24868\
        );

    \I__5571\ : InMux
    port map (
            O => \N__24890\,
            I => \N__24865\
        );

    \I__5570\ : InMux
    port map (
            O => \N__24889\,
            I => \N__24856\
        );

    \I__5569\ : InMux
    port map (
            O => \N__24888\,
            I => \N__24856\
        );

    \I__5568\ : InMux
    port map (
            O => \N__24887\,
            I => \N__24849\
        );

    \I__5567\ : InMux
    port map (
            O => \N__24886\,
            I => \N__24849\
        );

    \I__5566\ : InMux
    port map (
            O => \N__24885\,
            I => \N__24849\
        );

    \I__5565\ : InMux
    port map (
            O => \N__24882\,
            I => \N__24844\
        );

    \I__5564\ : InMux
    port map (
            O => \N__24879\,
            I => \N__24844\
        );

    \I__5563\ : InMux
    port map (
            O => \N__24878\,
            I => \N__24841\
        );

    \I__5562\ : InMux
    port map (
            O => \N__24875\,
            I => \N__24838\
        );

    \I__5561\ : InMux
    port map (
            O => \N__24874\,
            I => \N__24835\
        );

    \I__5560\ : LocalMux
    port map (
            O => \N__24871\,
            I => \N__24830\
        );

    \I__5559\ : LocalMux
    port map (
            O => \N__24868\,
            I => \N__24830\
        );

    \I__5558\ : LocalMux
    port map (
            O => \N__24865\,
            I => \N__24827\
        );

    \I__5557\ : InMux
    port map (
            O => \N__24864\,
            I => \N__24824\
        );

    \I__5556\ : InMux
    port map (
            O => \N__24863\,
            I => \N__24819\
        );

    \I__5555\ : InMux
    port map (
            O => \N__24862\,
            I => \N__24819\
        );

    \I__5554\ : CascadeMux
    port map (
            O => \N__24861\,
            I => \N__24816\
        );

    \I__5553\ : LocalMux
    port map (
            O => \N__24856\,
            I => \N__24810\
        );

    \I__5552\ : LocalMux
    port map (
            O => \N__24849\,
            I => \N__24807\
        );

    \I__5551\ : LocalMux
    port map (
            O => \N__24844\,
            I => \N__24804\
        );

    \I__5550\ : LocalMux
    port map (
            O => \N__24841\,
            I => \N__24797\
        );

    \I__5549\ : LocalMux
    port map (
            O => \N__24838\,
            I => \N__24797\
        );

    \I__5548\ : LocalMux
    port map (
            O => \N__24835\,
            I => \N__24790\
        );

    \I__5547\ : Span4Mux_s3_h
    port map (
            O => \N__24830\,
            I => \N__24790\
        );

    \I__5546\ : Span4Mux_h
    port map (
            O => \N__24827\,
            I => \N__24790\
        );

    \I__5545\ : LocalMux
    port map (
            O => \N__24824\,
            I => \N__24787\
        );

    \I__5544\ : LocalMux
    port map (
            O => \N__24819\,
            I => \N__24784\
        );

    \I__5543\ : InMux
    port map (
            O => \N__24816\,
            I => \N__24779\
        );

    \I__5542\ : InMux
    port map (
            O => \N__24815\,
            I => \N__24779\
        );

    \I__5541\ : InMux
    port map (
            O => \N__24814\,
            I => \N__24774\
        );

    \I__5540\ : InMux
    port map (
            O => \N__24813\,
            I => \N__24774\
        );

    \I__5539\ : Span4Mux_v
    port map (
            O => \N__24810\,
            I => \N__24767\
        );

    \I__5538\ : Span4Mux_h
    port map (
            O => \N__24807\,
            I => \N__24767\
        );

    \I__5537\ : Span4Mux_v
    port map (
            O => \N__24804\,
            I => \N__24767\
        );

    \I__5536\ : InMux
    port map (
            O => \N__24803\,
            I => \N__24762\
        );

    \I__5535\ : InMux
    port map (
            O => \N__24802\,
            I => \N__24762\
        );

    \I__5534\ : Span4Mux_s3_h
    port map (
            O => \N__24797\,
            I => \N__24757\
        );

    \I__5533\ : Span4Mux_h
    port map (
            O => \N__24790\,
            I => \N__24757\
        );

    \I__5532\ : Odrv4
    port map (
            O => \N__24787\,
            I => \Lab_UT.dictrl.currState_i_5_3\
        );

    \I__5531\ : Odrv4
    port map (
            O => \N__24784\,
            I => \Lab_UT.dictrl.currState_i_5_3\
        );

    \I__5530\ : LocalMux
    port map (
            O => \N__24779\,
            I => \Lab_UT.dictrl.currState_i_5_3\
        );

    \I__5529\ : LocalMux
    port map (
            O => \N__24774\,
            I => \Lab_UT.dictrl.currState_i_5_3\
        );

    \I__5528\ : Odrv4
    port map (
            O => \N__24767\,
            I => \Lab_UT.dictrl.currState_i_5_3\
        );

    \I__5527\ : LocalMux
    port map (
            O => \N__24762\,
            I => \Lab_UT.dictrl.currState_i_5_3\
        );

    \I__5526\ : Odrv4
    port map (
            O => \N__24757\,
            I => \Lab_UT.dictrl.currState_i_5_3\
        );

    \I__5525\ : CascadeMux
    port map (
            O => \N__24742\,
            I => \N__24739\
        );

    \I__5524\ : InMux
    port map (
            O => \N__24739\,
            I => \N__24736\
        );

    \I__5523\ : LocalMux
    port map (
            O => \N__24736\,
            I => \N__24733\
        );

    \I__5522\ : Odrv4
    port map (
            O => \N__24733\,
            I => \Lab_UT.dictrl.r_dicRun_r_1\
        );

    \I__5521\ : CascadeMux
    port map (
            O => \N__24730\,
            I => \N__24727\
        );

    \I__5520\ : InMux
    port map (
            O => \N__24727\,
            I => \N__24720\
        );

    \I__5519\ : InMux
    port map (
            O => \N__24726\,
            I => \N__24720\
        );

    \I__5518\ : InMux
    port map (
            O => \N__24725\,
            I => \N__24717\
        );

    \I__5517\ : LocalMux
    port map (
            O => \N__24720\,
            I => \N__24714\
        );

    \I__5516\ : LocalMux
    port map (
            O => \N__24717\,
            I => \N__24711\
        );

    \I__5515\ : Odrv4
    port map (
            O => \N__24714\,
            I => \Lab_UT.dictrl.r_dicLdMtens15_1i\
        );

    \I__5514\ : Odrv4
    port map (
            O => \N__24711\,
            I => \Lab_UT.dictrl.r_dicLdMtens15_1i\
        );

    \I__5513\ : InMux
    port map (
            O => \N__24706\,
            I => \N__24699\
        );

    \I__5512\ : InMux
    port map (
            O => \N__24705\,
            I => \N__24696\
        );

    \I__5511\ : InMux
    port map (
            O => \N__24704\,
            I => \N__24690\
        );

    \I__5510\ : InMux
    port map (
            O => \N__24703\,
            I => \N__24690\
        );

    \I__5509\ : IoInMux
    port map (
            O => \N__24702\,
            I => \N__24666\
        );

    \I__5508\ : LocalMux
    port map (
            O => \N__24699\,
            I => \N__24663\
        );

    \I__5507\ : LocalMux
    port map (
            O => \N__24696\,
            I => \N__24660\
        );

    \I__5506\ : InMux
    port map (
            O => \N__24695\,
            I => \N__24657\
        );

    \I__5505\ : LocalMux
    port map (
            O => \N__24690\,
            I => \N__24654\
        );

    \I__5504\ : InMux
    port map (
            O => \N__24689\,
            I => \N__24651\
        );

    \I__5503\ : InMux
    port map (
            O => \N__24688\,
            I => \N__24644\
        );

    \I__5502\ : InMux
    port map (
            O => \N__24687\,
            I => \N__24644\
        );

    \I__5501\ : InMux
    port map (
            O => \N__24686\,
            I => \N__24644\
        );

    \I__5500\ : InMux
    port map (
            O => \N__24685\,
            I => \N__24637\
        );

    \I__5499\ : InMux
    port map (
            O => \N__24684\,
            I => \N__24637\
        );

    \I__5498\ : InMux
    port map (
            O => \N__24683\,
            I => \N__24637\
        );

    \I__5497\ : InMux
    port map (
            O => \N__24682\,
            I => \N__24634\
        );

    \I__5496\ : InMux
    port map (
            O => \N__24681\,
            I => \N__24631\
        );

    \I__5495\ : InMux
    port map (
            O => \N__24680\,
            I => \N__24628\
        );

    \I__5494\ : InMux
    port map (
            O => \N__24679\,
            I => \N__24623\
        );

    \I__5493\ : InMux
    port map (
            O => \N__24678\,
            I => \N__24618\
        );

    \I__5492\ : InMux
    port map (
            O => \N__24677\,
            I => \N__24618\
        );

    \I__5491\ : InMux
    port map (
            O => \N__24676\,
            I => \N__24615\
        );

    \I__5490\ : InMux
    port map (
            O => \N__24675\,
            I => \N__24606\
        );

    \I__5489\ : InMux
    port map (
            O => \N__24674\,
            I => \N__24606\
        );

    \I__5488\ : InMux
    port map (
            O => \N__24673\,
            I => \N__24606\
        );

    \I__5487\ : InMux
    port map (
            O => \N__24672\,
            I => \N__24606\
        );

    \I__5486\ : InMux
    port map (
            O => \N__24671\,
            I => \N__24599\
        );

    \I__5485\ : InMux
    port map (
            O => \N__24670\,
            I => \N__24599\
        );

    \I__5484\ : InMux
    port map (
            O => \N__24669\,
            I => \N__24599\
        );

    \I__5483\ : LocalMux
    port map (
            O => \N__24666\,
            I => \N__24596\
        );

    \I__5482\ : Span4Mux_v
    port map (
            O => \N__24663\,
            I => \N__24591\
        );

    \I__5481\ : Span4Mux_v
    port map (
            O => \N__24660\,
            I => \N__24591\
        );

    \I__5480\ : LocalMux
    port map (
            O => \N__24657\,
            I => \N__24584\
        );

    \I__5479\ : Span4Mux_s3_v
    port map (
            O => \N__24654\,
            I => \N__24584\
        );

    \I__5478\ : LocalMux
    port map (
            O => \N__24651\,
            I => \N__24584\
        );

    \I__5477\ : LocalMux
    port map (
            O => \N__24644\,
            I => \N__24579\
        );

    \I__5476\ : LocalMux
    port map (
            O => \N__24637\,
            I => \N__24579\
        );

    \I__5475\ : LocalMux
    port map (
            O => \N__24634\,
            I => \N__24574\
        );

    \I__5474\ : LocalMux
    port map (
            O => \N__24631\,
            I => \N__24569\
        );

    \I__5473\ : LocalMux
    port map (
            O => \N__24628\,
            I => \N__24569\
        );

    \I__5472\ : InMux
    port map (
            O => \N__24627\,
            I => \N__24564\
        );

    \I__5471\ : InMux
    port map (
            O => \N__24626\,
            I => \N__24564\
        );

    \I__5470\ : LocalMux
    port map (
            O => \N__24623\,
            I => \N__24557\
        );

    \I__5469\ : LocalMux
    port map (
            O => \N__24618\,
            I => \N__24557\
        );

    \I__5468\ : LocalMux
    port map (
            O => \N__24615\,
            I => \N__24557\
        );

    \I__5467\ : LocalMux
    port map (
            O => \N__24606\,
            I => \N__24550\
        );

    \I__5466\ : LocalMux
    port map (
            O => \N__24599\,
            I => \N__24550\
        );

    \I__5465\ : IoSpan4Mux
    port map (
            O => \N__24596\,
            I => \N__24550\
        );

    \I__5464\ : Span4Mux_h
    port map (
            O => \N__24591\,
            I => \N__24547\
        );

    \I__5463\ : Span4Mux_v
    port map (
            O => \N__24584\,
            I => \N__24542\
        );

    \I__5462\ : Span4Mux_v
    port map (
            O => \N__24579\,
            I => \N__24542\
        );

    \I__5461\ : InMux
    port map (
            O => \N__24578\,
            I => \N__24537\
        );

    \I__5460\ : InMux
    port map (
            O => \N__24577\,
            I => \N__24537\
        );

    \I__5459\ : Span4Mux_h
    port map (
            O => \N__24574\,
            I => \N__24532\
        );

    \I__5458\ : Span4Mux_s3_h
    port map (
            O => \N__24569\,
            I => \N__24532\
        );

    \I__5457\ : LocalMux
    port map (
            O => \N__24564\,
            I => \N__24525\
        );

    \I__5456\ : Span4Mux_h
    port map (
            O => \N__24557\,
            I => \N__24525\
        );

    \I__5455\ : Span4Mux_s3_h
    port map (
            O => \N__24550\,
            I => \N__24525\
        );

    \I__5454\ : Odrv4
    port map (
            O => \N__24547\,
            I => rst
        );

    \I__5453\ : Odrv4
    port map (
            O => \N__24542\,
            I => rst
        );

    \I__5452\ : LocalMux
    port map (
            O => \N__24537\,
            I => rst
        );

    \I__5451\ : Odrv4
    port map (
            O => \N__24532\,
            I => rst
        );

    \I__5450\ : Odrv4
    port map (
            O => \N__24525\,
            I => rst
        );

    \I__5449\ : InMux
    port map (
            O => \N__24514\,
            I => \N__24509\
        );

    \I__5448\ : InMux
    port map (
            O => \N__24513\,
            I => \N__24504\
        );

    \I__5447\ : InMux
    port map (
            O => \N__24512\,
            I => \N__24504\
        );

    \I__5446\ : LocalMux
    port map (
            O => \N__24509\,
            I => \Lab_UT.dictrl.r_dicLdMtens15_1\
        );

    \I__5445\ : LocalMux
    port map (
            O => \N__24504\,
            I => \Lab_UT.dictrl.r_dicLdMtens15_1\
        );

    \I__5444\ : CascadeMux
    port map (
            O => \N__24499\,
            I => \Lab_UT.dictrl.decoder.de_atSignZ0Z_4_cascade_\
        );

    \I__5443\ : InMux
    port map (
            O => \N__24496\,
            I => \N__24490\
        );

    \I__5442\ : InMux
    port map (
            O => \N__24495\,
            I => \N__24490\
        );

    \I__5441\ : LocalMux
    port map (
            O => \N__24490\,
            I => \N__24487\
        );

    \I__5440\ : Odrv4
    port map (
            O => \N__24487\,
            I => \Lab_UT.dictrl.de_atSign\
        );

    \I__5439\ : CascadeMux
    port map (
            O => \N__24484\,
            I => \Lab_UT.dictrl.de_littleA_2_cascade_\
        );

    \I__5438\ : InMux
    port map (
            O => \N__24481\,
            I => \N__24478\
        );

    \I__5437\ : LocalMux
    port map (
            O => \N__24478\,
            I => \N__24472\
        );

    \I__5436\ : InMux
    port map (
            O => \N__24477\,
            I => \N__24469\
        );

    \I__5435\ : InMux
    port map (
            O => \N__24476\,
            I => \N__24466\
        );

    \I__5434\ : InMux
    port map (
            O => \N__24475\,
            I => \N__24463\
        );

    \I__5433\ : Span4Mux_h
    port map (
            O => \N__24472\,
            I => \N__24460\
        );

    \I__5432\ : LocalMux
    port map (
            O => \N__24469\,
            I => \N__24457\
        );

    \I__5431\ : LocalMux
    port map (
            O => \N__24466\,
            I => \Lab_UT.dictrl.de_littleL\
        );

    \I__5430\ : LocalMux
    port map (
            O => \N__24463\,
            I => \Lab_UT.dictrl.de_littleL\
        );

    \I__5429\ : Odrv4
    port map (
            O => \N__24460\,
            I => \Lab_UT.dictrl.de_littleL\
        );

    \I__5428\ : Odrv12
    port map (
            O => \N__24457\,
            I => \Lab_UT.dictrl.de_littleL\
        );

    \I__5427\ : InMux
    port map (
            O => \N__24448\,
            I => \N__24437\
        );

    \I__5426\ : InMux
    port map (
            O => \N__24447\,
            I => \N__24434\
        );

    \I__5425\ : InMux
    port map (
            O => \N__24446\,
            I => \N__24429\
        );

    \I__5424\ : InMux
    port map (
            O => \N__24445\,
            I => \N__24429\
        );

    \I__5423\ : InMux
    port map (
            O => \N__24444\,
            I => \N__24426\
        );

    \I__5422\ : InMux
    port map (
            O => \N__24443\,
            I => \N__24423\
        );

    \I__5421\ : InMux
    port map (
            O => \N__24442\,
            I => \N__24418\
        );

    \I__5420\ : InMux
    port map (
            O => \N__24441\,
            I => \N__24418\
        );

    \I__5419\ : InMux
    port map (
            O => \N__24440\,
            I => \N__24411\
        );

    \I__5418\ : LocalMux
    port map (
            O => \N__24437\,
            I => \N__24408\
        );

    \I__5417\ : LocalMux
    port map (
            O => \N__24434\,
            I => \N__24401\
        );

    \I__5416\ : LocalMux
    port map (
            O => \N__24429\,
            I => \N__24401\
        );

    \I__5415\ : LocalMux
    port map (
            O => \N__24426\,
            I => \N__24401\
        );

    \I__5414\ : LocalMux
    port map (
            O => \N__24423\,
            I => \N__24398\
        );

    \I__5413\ : LocalMux
    port map (
            O => \N__24418\,
            I => \N__24395\
        );

    \I__5412\ : InMux
    port map (
            O => \N__24417\,
            I => \N__24392\
        );

    \I__5411\ : InMux
    port map (
            O => \N__24416\,
            I => \N__24387\
        );

    \I__5410\ : InMux
    port map (
            O => \N__24415\,
            I => \N__24387\
        );

    \I__5409\ : InMux
    port map (
            O => \N__24414\,
            I => \N__24384\
        );

    \I__5408\ : LocalMux
    port map (
            O => \N__24411\,
            I => \N__24379\
        );

    \I__5407\ : Span4Mux_v
    port map (
            O => \N__24408\,
            I => \N__24379\
        );

    \I__5406\ : Span4Mux_h
    port map (
            O => \N__24401\,
            I => \N__24376\
        );

    \I__5405\ : Span4Mux_h
    port map (
            O => \N__24398\,
            I => \N__24371\
        );

    \I__5404\ : Span4Mux_s2_v
    port map (
            O => \N__24395\,
            I => \N__24371\
        );

    \I__5403\ : LocalMux
    port map (
            O => \N__24392\,
            I => bu_rx_data_5
        );

    \I__5402\ : LocalMux
    port map (
            O => \N__24387\,
            I => bu_rx_data_5
        );

    \I__5401\ : LocalMux
    port map (
            O => \N__24384\,
            I => bu_rx_data_5
        );

    \I__5400\ : Odrv4
    port map (
            O => \N__24379\,
            I => bu_rx_data_5
        );

    \I__5399\ : Odrv4
    port map (
            O => \N__24376\,
            I => bu_rx_data_5
        );

    \I__5398\ : Odrv4
    port map (
            O => \N__24371\,
            I => bu_rx_data_5
        );

    \I__5397\ : InMux
    port map (
            O => \N__24358\,
            I => \N__24351\
        );

    \I__5396\ : InMux
    port map (
            O => \N__24357\,
            I => \N__24351\
        );

    \I__5395\ : InMux
    port map (
            O => \N__24356\,
            I => \N__24348\
        );

    \I__5394\ : LocalMux
    port map (
            O => \N__24351\,
            I => \N__24344\
        );

    \I__5393\ : LocalMux
    port map (
            O => \N__24348\,
            I => \N__24341\
        );

    \I__5392\ : InMux
    port map (
            O => \N__24347\,
            I => \N__24337\
        );

    \I__5391\ : Span4Mux_v
    port map (
            O => \N__24344\,
            I => \N__24332\
        );

    \I__5390\ : Span4Mux_s2_v
    port map (
            O => \N__24341\,
            I => \N__24332\
        );

    \I__5389\ : InMux
    port map (
            O => \N__24340\,
            I => \N__24329\
        );

    \I__5388\ : LocalMux
    port map (
            O => \N__24337\,
            I => \Lab_UT.dictrl.de_littleL_4\
        );

    \I__5387\ : Odrv4
    port map (
            O => \N__24332\,
            I => \Lab_UT.dictrl.de_littleL_4\
        );

    \I__5386\ : LocalMux
    port map (
            O => \N__24329\,
            I => \Lab_UT.dictrl.de_littleL_4\
        );

    \I__5385\ : CascadeMux
    port map (
            O => \N__24322\,
            I => \N__24317\
        );

    \I__5384\ : CascadeMux
    port map (
            O => \N__24321\,
            I => \N__24314\
        );

    \I__5383\ : CascadeMux
    port map (
            O => \N__24320\,
            I => \N__24311\
        );

    \I__5382\ : InMux
    port map (
            O => \N__24317\,
            I => \N__24301\
        );

    \I__5381\ : InMux
    port map (
            O => \N__24314\,
            I => \N__24301\
        );

    \I__5380\ : InMux
    port map (
            O => \N__24311\,
            I => \N__24301\
        );

    \I__5379\ : CascadeMux
    port map (
            O => \N__24310\,
            I => \N__24297\
        );

    \I__5378\ : InMux
    port map (
            O => \N__24309\,
            I => \N__24291\
        );

    \I__5377\ : InMux
    port map (
            O => \N__24308\,
            I => \N__24288\
        );

    \I__5376\ : LocalMux
    port map (
            O => \N__24301\,
            I => \N__24285\
        );

    \I__5375\ : InMux
    port map (
            O => \N__24300\,
            I => \N__24282\
        );

    \I__5374\ : InMux
    port map (
            O => \N__24297\,
            I => \N__24275\
        );

    \I__5373\ : InMux
    port map (
            O => \N__24296\,
            I => \N__24275\
        );

    \I__5372\ : InMux
    port map (
            O => \N__24295\,
            I => \N__24275\
        );

    \I__5371\ : CascadeMux
    port map (
            O => \N__24294\,
            I => \N__24272\
        );

    \I__5370\ : LocalMux
    port map (
            O => \N__24291\,
            I => \N__24267\
        );

    \I__5369\ : LocalMux
    port map (
            O => \N__24288\,
            I => \N__24263\
        );

    \I__5368\ : Span4Mux_s3_h
    port map (
            O => \N__24285\,
            I => \N__24260\
        );

    \I__5367\ : LocalMux
    port map (
            O => \N__24282\,
            I => \N__24255\
        );

    \I__5366\ : LocalMux
    port map (
            O => \N__24275\,
            I => \N__24255\
        );

    \I__5365\ : InMux
    port map (
            O => \N__24272\,
            I => \N__24252\
        );

    \I__5364\ : InMux
    port map (
            O => \N__24271\,
            I => \N__24247\
        );

    \I__5363\ : InMux
    port map (
            O => \N__24270\,
            I => \N__24247\
        );

    \I__5362\ : Span4Mux_v
    port map (
            O => \N__24267\,
            I => \N__24244\
        );

    \I__5361\ : InMux
    port map (
            O => \N__24266\,
            I => \N__24241\
        );

    \I__5360\ : Span4Mux_h
    port map (
            O => \N__24263\,
            I => \N__24238\
        );

    \I__5359\ : Span4Mux_h
    port map (
            O => \N__24260\,
            I => \N__24235\
        );

    \I__5358\ : Span4Mux_v
    port map (
            O => \N__24255\,
            I => \N__24230\
        );

    \I__5357\ : LocalMux
    port map (
            O => \N__24252\,
            I => \N__24230\
        );

    \I__5356\ : LocalMux
    port map (
            O => \N__24247\,
            I => bu_rx_data_6
        );

    \I__5355\ : Odrv4
    port map (
            O => \N__24244\,
            I => bu_rx_data_6
        );

    \I__5354\ : LocalMux
    port map (
            O => \N__24241\,
            I => bu_rx_data_6
        );

    \I__5353\ : Odrv4
    port map (
            O => \N__24238\,
            I => bu_rx_data_6
        );

    \I__5352\ : Odrv4
    port map (
            O => \N__24235\,
            I => bu_rx_data_6
        );

    \I__5351\ : Odrv4
    port map (
            O => \N__24230\,
            I => bu_rx_data_6
        );

    \I__5350\ : InMux
    port map (
            O => \N__24217\,
            I => \N__24214\
        );

    \I__5349\ : LocalMux
    port map (
            O => \N__24214\,
            I => \N__24211\
        );

    \I__5348\ : Odrv4
    port map (
            O => \N__24211\,
            I => \Lab_UT.dictrl.g0_4_2\
        );

    \I__5347\ : CascadeMux
    port map (
            O => \N__24208\,
            I => \N__24203\
        );

    \I__5346\ : InMux
    port map (
            O => \N__24207\,
            I => \N__24200\
        );

    \I__5345\ : CascadeMux
    port map (
            O => \N__24206\,
            I => \N__24197\
        );

    \I__5344\ : InMux
    port map (
            O => \N__24203\,
            I => \N__24194\
        );

    \I__5343\ : LocalMux
    port map (
            O => \N__24200\,
            I => \N__24191\
        );

    \I__5342\ : InMux
    port map (
            O => \N__24197\,
            I => \N__24188\
        );

    \I__5341\ : LocalMux
    port map (
            O => \N__24194\,
            I => \N__24185\
        );

    \I__5340\ : Odrv12
    port map (
            O => \N__24191\,
            I => \Lab_UT.dictrl.de_littleA_2\
        );

    \I__5339\ : LocalMux
    port map (
            O => \N__24188\,
            I => \Lab_UT.dictrl.de_littleA_2\
        );

    \I__5338\ : Odrv4
    port map (
            O => \N__24185\,
            I => \Lab_UT.dictrl.de_littleA_2\
        );

    \I__5337\ : InMux
    port map (
            O => \N__24178\,
            I => \N__24173\
        );

    \I__5336\ : CascadeMux
    port map (
            O => \N__24177\,
            I => \N__24169\
        );

    \I__5335\ : CascadeMux
    port map (
            O => \N__24176\,
            I => \N__24165\
        );

    \I__5334\ : LocalMux
    port map (
            O => \N__24173\,
            I => \N__24162\
        );

    \I__5333\ : InMux
    port map (
            O => \N__24172\,
            I => \N__24159\
        );

    \I__5332\ : InMux
    port map (
            O => \N__24169\,
            I => \N__24150\
        );

    \I__5331\ : InMux
    port map (
            O => \N__24168\,
            I => \N__24150\
        );

    \I__5330\ : InMux
    port map (
            O => \N__24165\,
            I => \N__24150\
        );

    \I__5329\ : Span4Mux_h
    port map (
            O => \N__24162\,
            I => \N__24145\
        );

    \I__5328\ : LocalMux
    port map (
            O => \N__24159\,
            I => \N__24145\
        );

    \I__5327\ : InMux
    port map (
            O => \N__24158\,
            I => \N__24140\
        );

    \I__5326\ : InMux
    port map (
            O => \N__24157\,
            I => \N__24140\
        );

    \I__5325\ : LocalMux
    port map (
            O => \N__24150\,
            I => \Lab_UT.dictrl.un2_dicAlarmTrig\
        );

    \I__5324\ : Odrv4
    port map (
            O => \N__24145\,
            I => \Lab_UT.dictrl.un2_dicAlarmTrig\
        );

    \I__5323\ : LocalMux
    port map (
            O => \N__24140\,
            I => \Lab_UT.dictrl.un2_dicAlarmTrig\
        );

    \I__5322\ : InMux
    port map (
            O => \N__24133\,
            I => \N__24130\
        );

    \I__5321\ : LocalMux
    port map (
            O => \N__24130\,
            I => \Lab_UT.dictrl.N_186\
        );

    \I__5320\ : CascadeMux
    port map (
            O => \N__24127\,
            I => \N__24123\
        );

    \I__5319\ : InMux
    port map (
            O => \N__24126\,
            I => \N__24113\
        );

    \I__5318\ : InMux
    port map (
            O => \N__24123\,
            I => \N__24113\
        );

    \I__5317\ : InMux
    port map (
            O => \N__24122\,
            I => \N__24113\
        );

    \I__5316\ : CascadeMux
    port map (
            O => \N__24121\,
            I => \N__24110\
        );

    \I__5315\ : CascadeMux
    port map (
            O => \N__24120\,
            I => \N__24107\
        );

    \I__5314\ : LocalMux
    port map (
            O => \N__24113\,
            I => \N__24104\
        );

    \I__5313\ : InMux
    port map (
            O => \N__24110\,
            I => \N__24101\
        );

    \I__5312\ : InMux
    port map (
            O => \N__24107\,
            I => \N__24098\
        );

    \I__5311\ : Span4Mux_h
    port map (
            O => \N__24104\,
            I => \N__24095\
        );

    \I__5310\ : LocalMux
    port map (
            O => \N__24101\,
            I => \Lab_UT.dictrl.nextState_al_0_0\
        );

    \I__5309\ : LocalMux
    port map (
            O => \N__24098\,
            I => \Lab_UT.dictrl.nextState_al_0_0\
        );

    \I__5308\ : Odrv4
    port map (
            O => \N__24095\,
            I => \Lab_UT.dictrl.nextState_al_0_0\
        );

    \I__5307\ : CascadeMux
    port map (
            O => \N__24088\,
            I => \Lab_UT.dictrl.N_186_cascade_\
        );

    \I__5306\ : InMux
    port map (
            O => \N__24085\,
            I => \N__24081\
        );

    \I__5305\ : InMux
    port map (
            O => \N__24084\,
            I => \N__24078\
        );

    \I__5304\ : LocalMux
    port map (
            O => \N__24081\,
            I => \Lab_UT.dictrl.nextState_al_1_0_0_1\
        );

    \I__5303\ : LocalMux
    port map (
            O => \N__24078\,
            I => \Lab_UT.dictrl.nextState_al_1_0_0_1\
        );

    \I__5302\ : CascadeMux
    port map (
            O => \N__24073\,
            I => \N__24069\
        );

    \I__5301\ : InMux
    port map (
            O => \N__24072\,
            I => \N__24061\
        );

    \I__5300\ : InMux
    port map (
            O => \N__24069\,
            I => \N__24061\
        );

    \I__5299\ : InMux
    port map (
            O => \N__24068\,
            I => \N__24061\
        );

    \I__5298\ : LocalMux
    port map (
            O => \N__24061\,
            I => \Lab_UT.dictrl.currState_alZ0Z_0\
        );

    \I__5297\ : InMux
    port map (
            O => \N__24058\,
            I => \N__24047\
        );

    \I__5296\ : InMux
    port map (
            O => \N__24057\,
            I => \N__24047\
        );

    \I__5295\ : InMux
    port map (
            O => \N__24056\,
            I => \N__24044\
        );

    \I__5294\ : InMux
    port map (
            O => \N__24055\,
            I => \N__24035\
        );

    \I__5293\ : InMux
    port map (
            O => \N__24054\,
            I => \N__24035\
        );

    \I__5292\ : InMux
    port map (
            O => \N__24053\,
            I => \N__24035\
        );

    \I__5291\ : InMux
    port map (
            O => \N__24052\,
            I => \N__24035\
        );

    \I__5290\ : LocalMux
    port map (
            O => \N__24047\,
            I => \Lab_UT.dictrl.currState_alZ0Z_1\
        );

    \I__5289\ : LocalMux
    port map (
            O => \N__24044\,
            I => \Lab_UT.dictrl.currState_alZ0Z_1\
        );

    \I__5288\ : LocalMux
    port map (
            O => \N__24035\,
            I => \Lab_UT.dictrl.currState_alZ0Z_1\
        );

    \I__5287\ : CascadeMux
    port map (
            O => \N__24028\,
            I => \N__24025\
        );

    \I__5286\ : InMux
    port map (
            O => \N__24025\,
            I => \N__24022\
        );

    \I__5285\ : LocalMux
    port map (
            O => \N__24022\,
            I => \N__24019\
        );

    \I__5284\ : Span12Mux_s11_h
    port map (
            O => \N__24019\,
            I => \N__24016\
        );

    \I__5283\ : Odrv12
    port map (
            O => \N__24016\,
            I => \Lab_UT.dictrl.currState_i_5_1\
        );

    \I__5282\ : InMux
    port map (
            O => \N__24013\,
            I => \N__24008\
        );

    \I__5281\ : CascadeMux
    port map (
            O => \N__24012\,
            I => \N__24000\
        );

    \I__5280\ : InMux
    port map (
            O => \N__24011\,
            I => \N__23997\
        );

    \I__5279\ : LocalMux
    port map (
            O => \N__24008\,
            I => \N__23994\
        );

    \I__5278\ : InMux
    port map (
            O => \N__24007\,
            I => \N__23991\
        );

    \I__5277\ : InMux
    port map (
            O => \N__24006\,
            I => \N__23988\
        );

    \I__5276\ : InMux
    port map (
            O => \N__24005\,
            I => \N__23985\
        );

    \I__5275\ : InMux
    port map (
            O => \N__24004\,
            I => \N__23982\
        );

    \I__5274\ : InMux
    port map (
            O => \N__24003\,
            I => \N__23977\
        );

    \I__5273\ : InMux
    port map (
            O => \N__24000\,
            I => \N__23977\
        );

    \I__5272\ : LocalMux
    port map (
            O => \N__23997\,
            I => \N__23973\
        );

    \I__5271\ : Span4Mux_v
    port map (
            O => \N__23994\,
            I => \N__23969\
        );

    \I__5270\ : LocalMux
    port map (
            O => \N__23991\,
            I => \N__23966\
        );

    \I__5269\ : LocalMux
    port map (
            O => \N__23988\,
            I => \N__23963\
        );

    \I__5268\ : LocalMux
    port map (
            O => \N__23985\,
            I => \N__23960\
        );

    \I__5267\ : LocalMux
    port map (
            O => \N__23982\,
            I => \N__23955\
        );

    \I__5266\ : LocalMux
    port map (
            O => \N__23977\,
            I => \N__23955\
        );

    \I__5265\ : InMux
    port map (
            O => \N__23976\,
            I => \N__23952\
        );

    \I__5264\ : Span4Mux_v
    port map (
            O => \N__23973\,
            I => \N__23949\
        );

    \I__5263\ : InMux
    port map (
            O => \N__23972\,
            I => \N__23946\
        );

    \I__5262\ : Span4Mux_h
    port map (
            O => \N__23969\,
            I => \N__23937\
        );

    \I__5261\ : Span4Mux_v
    port map (
            O => \N__23966\,
            I => \N__23937\
        );

    \I__5260\ : Span4Mux_v
    port map (
            O => \N__23963\,
            I => \N__23937\
        );

    \I__5259\ : Span4Mux_v
    port map (
            O => \N__23960\,
            I => \N__23937\
        );

    \I__5258\ : Span4Mux_v
    port map (
            O => \N__23955\,
            I => \N__23934\
        );

    \I__5257\ : LocalMux
    port map (
            O => \N__23952\,
            I => \Lab_UT.dictrl.currState_i_5_0\
        );

    \I__5256\ : Odrv4
    port map (
            O => \N__23949\,
            I => \Lab_UT.dictrl.currState_i_5_0\
        );

    \I__5255\ : LocalMux
    port map (
            O => \N__23946\,
            I => \Lab_UT.dictrl.currState_i_5_0\
        );

    \I__5254\ : Odrv4
    port map (
            O => \N__23937\,
            I => \Lab_UT.dictrl.currState_i_5_0\
        );

    \I__5253\ : Odrv4
    port map (
            O => \N__23934\,
            I => \Lab_UT.dictrl.currState_i_5_0\
        );

    \I__5252\ : CascadeMux
    port map (
            O => \N__23923\,
            I => \Lab_UT.dictrl.un1_currState_8_u_ns_1_cascade_\
        );

    \I__5251\ : SRMux
    port map (
            O => \N__23920\,
            I => \N__23917\
        );

    \I__5250\ : LocalMux
    port map (
            O => \N__23917\,
            I => \N__23914\
        );

    \I__5249\ : Sp12to4
    port map (
            O => \N__23914\,
            I => \N__23910\
        );

    \I__5248\ : InMux
    port map (
            O => \N__23913\,
            I => \N__23907\
        );

    \I__5247\ : Odrv12
    port map (
            O => \N__23910\,
            I => \Lab_UT.dictrl.currState_ret_7_RNI03VHZ0Z1\
        );

    \I__5246\ : LocalMux
    port map (
            O => \N__23907\,
            I => \Lab_UT.dictrl.currState_ret_7_RNI03VHZ0Z1\
        );

    \I__5245\ : CascadeMux
    port map (
            O => \N__23902\,
            I => \Lab_UT.dictrl.un1_currState_inv_1_cascade_\
        );

    \I__5244\ : SRMux
    port map (
            O => \N__23899\,
            I => \N__23895\
        );

    \I__5243\ : InMux
    port map (
            O => \N__23898\,
            I => \N__23892\
        );

    \I__5242\ : LocalMux
    port map (
            O => \N__23895\,
            I => \N__23889\
        );

    \I__5241\ : LocalMux
    port map (
            O => \N__23892\,
            I => \N__23886\
        );

    \I__5240\ : Span4Mux_h
    port map (
            O => \N__23889\,
            I => \N__23883\
        );

    \I__5239\ : Span4Mux_v
    port map (
            O => \N__23886\,
            I => \N__23880\
        );

    \I__5238\ : Span4Mux_v
    port map (
            O => \N__23883\,
            I => \N__23877\
        );

    \I__5237\ : Span4Mux_h
    port map (
            O => \N__23880\,
            I => \N__23874\
        );

    \I__5236\ : Odrv4
    port map (
            O => \N__23877\,
            I => \Lab_UT.dictrl.currState_0_ret_1_RNIPH7FZ0Z1\
        );

    \I__5235\ : Odrv4
    port map (
            O => \N__23874\,
            I => \Lab_UT.dictrl.currState_0_ret_1_RNIPH7FZ0Z1\
        );

    \I__5234\ : InMux
    port map (
            O => \N__23869\,
            I => \N__23866\
        );

    \I__5233\ : LocalMux
    port map (
            O => \N__23866\,
            I => \N__23863\
        );

    \I__5232\ : Odrv12
    port map (
            O => \N__23863\,
            I => \Lab_UT.dictrl.r_dicLdMtens14_1\
        );

    \I__5231\ : InMux
    port map (
            O => \N__23860\,
            I => \N__23857\
        );

    \I__5230\ : LocalMux
    port map (
            O => \N__23857\,
            I => \N__23851\
        );

    \I__5229\ : InMux
    port map (
            O => \N__23856\,
            I => \N__23846\
        );

    \I__5228\ : InMux
    port map (
            O => \N__23855\,
            I => \N__23846\
        );

    \I__5227\ : InMux
    port map (
            O => \N__23854\,
            I => \N__23843\
        );

    \I__5226\ : Span4Mux_h
    port map (
            O => \N__23851\,
            I => \N__23836\
        );

    \I__5225\ : LocalMux
    port map (
            O => \N__23846\,
            I => \N__23836\
        );

    \I__5224\ : LocalMux
    port map (
            O => \N__23843\,
            I => \N__23836\
        );

    \I__5223\ : Odrv4
    port map (
            O => \N__23836\,
            I => \Lab_UT.dictrl.r_Sone_init5_1\
        );

    \I__5222\ : CascadeMux
    port map (
            O => \N__23833\,
            I => \N__23828\
        );

    \I__5221\ : InMux
    port map (
            O => \N__23832\,
            I => \N__23819\
        );

    \I__5220\ : InMux
    port map (
            O => \N__23831\,
            I => \N__23819\
        );

    \I__5219\ : InMux
    port map (
            O => \N__23828\,
            I => \N__23807\
        );

    \I__5218\ : InMux
    port map (
            O => \N__23827\,
            I => \N__23807\
        );

    \I__5217\ : InMux
    port map (
            O => \N__23826\,
            I => \N__23804\
        );

    \I__5216\ : InMux
    port map (
            O => \N__23825\,
            I => \N__23799\
        );

    \I__5215\ : InMux
    port map (
            O => \N__23824\,
            I => \N__23799\
        );

    \I__5214\ : LocalMux
    port map (
            O => \N__23819\,
            I => \N__23795\
        );

    \I__5213\ : InMux
    port map (
            O => \N__23818\,
            I => \N__23792\
        );

    \I__5212\ : InMux
    port map (
            O => \N__23817\,
            I => \N__23789\
        );

    \I__5211\ : InMux
    port map (
            O => \N__23816\,
            I => \N__23786\
        );

    \I__5210\ : InMux
    port map (
            O => \N__23815\,
            I => \N__23781\
        );

    \I__5209\ : InMux
    port map (
            O => \N__23814\,
            I => \N__23778\
        );

    \I__5208\ : InMux
    port map (
            O => \N__23813\,
            I => \N__23772\
        );

    \I__5207\ : InMux
    port map (
            O => \N__23812\,
            I => \N__23769\
        );

    \I__5206\ : LocalMux
    port map (
            O => \N__23807\,
            I => \N__23764\
        );

    \I__5205\ : LocalMux
    port map (
            O => \N__23804\,
            I => \N__23764\
        );

    \I__5204\ : LocalMux
    port map (
            O => \N__23799\,
            I => \N__23761\
        );

    \I__5203\ : InMux
    port map (
            O => \N__23798\,
            I => \N__23758\
        );

    \I__5202\ : Span4Mux_v
    port map (
            O => \N__23795\,
            I => \N__23749\
        );

    \I__5201\ : LocalMux
    port map (
            O => \N__23792\,
            I => \N__23749\
        );

    \I__5200\ : LocalMux
    port map (
            O => \N__23789\,
            I => \N__23749\
        );

    \I__5199\ : LocalMux
    port map (
            O => \N__23786\,
            I => \N__23749\
        );

    \I__5198\ : InMux
    port map (
            O => \N__23785\,
            I => \N__23744\
        );

    \I__5197\ : InMux
    port map (
            O => \N__23784\,
            I => \N__23744\
        );

    \I__5196\ : LocalMux
    port map (
            O => \N__23781\,
            I => \N__23741\
        );

    \I__5195\ : LocalMux
    port map (
            O => \N__23778\,
            I => \N__23738\
        );

    \I__5194\ : InMux
    port map (
            O => \N__23777\,
            I => \N__23731\
        );

    \I__5193\ : InMux
    port map (
            O => \N__23776\,
            I => \N__23731\
        );

    \I__5192\ : InMux
    port map (
            O => \N__23775\,
            I => \N__23731\
        );

    \I__5191\ : LocalMux
    port map (
            O => \N__23772\,
            I => \N__23724\
        );

    \I__5190\ : LocalMux
    port map (
            O => \N__23769\,
            I => \N__23724\
        );

    \I__5189\ : Span4Mux_h
    port map (
            O => \N__23764\,
            I => \N__23724\
        );

    \I__5188\ : Span4Mux_v
    port map (
            O => \N__23761\,
            I => \N__23721\
        );

    \I__5187\ : LocalMux
    port map (
            O => \N__23758\,
            I => \N__23716\
        );

    \I__5186\ : Span4Mux_h
    port map (
            O => \N__23749\,
            I => \N__23716\
        );

    \I__5185\ : LocalMux
    port map (
            O => \N__23744\,
            I => \N__23709\
        );

    \I__5184\ : Span4Mux_v
    port map (
            O => \N__23741\,
            I => \N__23709\
        );

    \I__5183\ : Span4Mux_s3_h
    port map (
            O => \N__23738\,
            I => \N__23709\
        );

    \I__5182\ : LocalMux
    port map (
            O => \N__23731\,
            I => \N__23704\
        );

    \I__5181\ : Span4Mux_h
    port map (
            O => \N__23724\,
            I => \N__23704\
        );

    \I__5180\ : Span4Mux_h
    port map (
            O => \N__23721\,
            I => \N__23699\
        );

    \I__5179\ : Span4Mux_v
    port map (
            O => \N__23716\,
            I => \N__23699\
        );

    \I__5178\ : Span4Mux_h
    port map (
            O => \N__23709\,
            I => \N__23696\
        );

    \I__5177\ : Span4Mux_v
    port map (
            O => \N__23704\,
            I => \N__23693\
        );

    \I__5176\ : Odrv4
    port map (
            O => \N__23699\,
            I => \Lab_UT.dictrl.currStateZ0Z_3\
        );

    \I__5175\ : Odrv4
    port map (
            O => \N__23696\,
            I => \Lab_UT.dictrl.currStateZ0Z_3\
        );

    \I__5174\ : Odrv4
    port map (
            O => \N__23693\,
            I => \Lab_UT.dictrl.currStateZ0Z_3\
        );

    \I__5173\ : InMux
    port map (
            O => \N__23686\,
            I => \N__23682\
        );

    \I__5172\ : InMux
    port map (
            O => \N__23685\,
            I => \N__23679\
        );

    \I__5171\ : LocalMux
    port map (
            O => \N__23682\,
            I => \Lab_UT.dictrl.un1_currState_inv_1\
        );

    \I__5170\ : LocalMux
    port map (
            O => \N__23679\,
            I => \Lab_UT.dictrl.un1_currState_inv_1\
        );

    \I__5169\ : CascadeMux
    port map (
            O => \N__23674\,
            I => \Lab_UT.dictrl.N_201_cascade_\
        );

    \I__5168\ : SRMux
    port map (
            O => \N__23671\,
            I => \N__23665\
        );

    \I__5167\ : InMux
    port map (
            O => \N__23670\,
            I => \N__23665\
        );

    \I__5166\ : LocalMux
    port map (
            O => \N__23665\,
            I => \N__23662\
        );

    \I__5165\ : Span4Mux_h
    port map (
            O => \N__23662\,
            I => \N__23659\
        );

    \I__5164\ : Odrv4
    port map (
            O => \N__23659\,
            I => \Lab_UT.dictrl.currState_2_RNIOB6H1Z0Z_2\
        );

    \I__5163\ : InMux
    port map (
            O => \N__23656\,
            I => \N__23647\
        );

    \I__5162\ : InMux
    port map (
            O => \N__23655\,
            I => \N__23647\
        );

    \I__5161\ : InMux
    port map (
            O => \N__23654\,
            I => \N__23647\
        );

    \I__5160\ : LocalMux
    port map (
            O => \N__23647\,
            I => \N__23642\
        );

    \I__5159\ : InMux
    port map (
            O => \N__23646\,
            I => \N__23639\
        );

    \I__5158\ : InMux
    port map (
            O => \N__23645\,
            I => \N__23634\
        );

    \I__5157\ : Span4Mux_h
    port map (
            O => \N__23642\,
            I => \N__23631\
        );

    \I__5156\ : LocalMux
    port map (
            O => \N__23639\,
            I => \N__23628\
        );

    \I__5155\ : InMux
    port map (
            O => \N__23638\,
            I => \N__23623\
        );

    \I__5154\ : InMux
    port map (
            O => \N__23637\,
            I => \N__23623\
        );

    \I__5153\ : LocalMux
    port map (
            O => \N__23634\,
            I => \Lab_UT.dictrl.r_dicAlarmTrigZ0\
        );

    \I__5152\ : Odrv4
    port map (
            O => \N__23631\,
            I => \Lab_UT.dictrl.r_dicAlarmTrigZ0\
        );

    \I__5151\ : Odrv4
    port map (
            O => \N__23628\,
            I => \Lab_UT.dictrl.r_dicAlarmTrigZ0\
        );

    \I__5150\ : LocalMux
    port map (
            O => \N__23623\,
            I => \Lab_UT.dictrl.r_dicAlarmTrigZ0\
        );

    \I__5149\ : InMux
    port map (
            O => \N__23614\,
            I => \N__23611\
        );

    \I__5148\ : LocalMux
    port map (
            O => \N__23611\,
            I => \N__23608\
        );

    \I__5147\ : Odrv12
    port map (
            O => \N__23608\,
            I => \Lab_UT.displayAlarmZ0Z_5\
        );

    \I__5146\ : InMux
    port map (
            O => \N__23605\,
            I => \N__23602\
        );

    \I__5145\ : LocalMux
    port map (
            O => \N__23602\,
            I => \Lab_UT.dictrl.nextState_al_1\
        );

    \I__5144\ : CascadeMux
    port map (
            O => \N__23599\,
            I => \Lab_UT.dictrl.nextState_al_1_cascade_\
        );

    \I__5143\ : CascadeMux
    port map (
            O => \N__23596\,
            I => \N__23592\
        );

    \I__5142\ : InMux
    port map (
            O => \N__23595\,
            I => \N__23589\
        );

    \I__5141\ : InMux
    port map (
            O => \N__23592\,
            I => \N__23586\
        );

    \I__5140\ : LocalMux
    port map (
            O => \N__23589\,
            I => \Lab_UT.dictrl.un2_dicAlarmTrig_i_6\
        );

    \I__5139\ : LocalMux
    port map (
            O => \N__23586\,
            I => \Lab_UT.dictrl.un2_dicAlarmTrig_i_6\
        );

    \I__5138\ : InMux
    port map (
            O => \N__23581\,
            I => \N__23578\
        );

    \I__5137\ : LocalMux
    port map (
            O => \N__23578\,
            I => \Lab_UT.dictrl.nextState_al_latmux_1\
        );

    \I__5136\ : CascadeMux
    port map (
            O => \N__23575\,
            I => \Lab_UT.dictrl.nextState_al_latmux_1_cascade_\
        );

    \I__5135\ : InMux
    port map (
            O => \N__23572\,
            I => \N__23566\
        );

    \I__5134\ : InMux
    port map (
            O => \N__23571\,
            I => \N__23566\
        );

    \I__5133\ : LocalMux
    port map (
            O => \N__23566\,
            I => \Lab_UT.dictrl.nextState_alZ0Z_0\
        );

    \I__5132\ : InMux
    port map (
            O => \N__23563\,
            I => \N__23560\
        );

    \I__5131\ : LocalMux
    port map (
            O => \N__23560\,
            I => \Lab_UT.didp.Stens_subtractor.un1_q_axb0\
        );

    \I__5130\ : InMux
    port map (
            O => \N__23557\,
            I => \N__23554\
        );

    \I__5129\ : LocalMux
    port map (
            O => \N__23554\,
            I => \Lab_UT.didp.Stens_subtractor.q_RNO_0_0_3\
        );

    \I__5128\ : InMux
    port map (
            O => \N__23551\,
            I => \N__23542\
        );

    \I__5127\ : InMux
    port map (
            O => \N__23550\,
            I => \N__23542\
        );

    \I__5126\ : InMux
    port map (
            O => \N__23549\,
            I => \N__23542\
        );

    \I__5125\ : LocalMux
    port map (
            O => \N__23542\,
            I => \Lab_UT.didp.Stens_subtractor.N_86\
        );

    \I__5124\ : InMux
    port map (
            O => \N__23539\,
            I => \N__23536\
        );

    \I__5123\ : LocalMux
    port map (
            O => \N__23536\,
            I => \Lab_UT.didp.Stens_subtractor.q_RNO_0_1_2\
        );

    \I__5122\ : CascadeMux
    port map (
            O => \N__23533\,
            I => \Lab_UT.didp.q_RNIDDF11_3_cascade_\
        );

    \I__5121\ : IoInMux
    port map (
            O => \N__23530\,
            I => \N__23527\
        );

    \I__5120\ : LocalMux
    port map (
            O => \N__23527\,
            I => \N__23524\
        );

    \I__5119\ : Span4Mux_s3_h
    port map (
            O => \N__23524\,
            I => \N__23521\
        );

    \I__5118\ : Odrv4
    port map (
            O => \N__23521\,
            I => led_c_3
        );

    \I__5117\ : InMux
    port map (
            O => \N__23518\,
            I => \N__23515\
        );

    \I__5116\ : LocalMux
    port map (
            O => \N__23515\,
            I => \Lab_UT.didp.q_RNI1TVP_3\
        );

    \I__5115\ : InMux
    port map (
            O => \N__23512\,
            I => \N__23509\
        );

    \I__5114\ : LocalMux
    port map (
            O => \N__23509\,
            I => \Lab_UT.didp.q_RNIBBF11_2\
        );

    \I__5113\ : InMux
    port map (
            O => \N__23506\,
            I => \N__23503\
        );

    \I__5112\ : LocalMux
    port map (
            O => \N__23503\,
            I => \N__23500\
        );

    \I__5111\ : Span4Mux_h
    port map (
            O => \N__23500\,
            I => \N__23497\
        );

    \I__5110\ : Odrv4
    port map (
            O => \N__23497\,
            I => \Lab_UT.didp.q_RNIVQVP_2\
        );

    \I__5109\ : IoInMux
    port map (
            O => \N__23494\,
            I => \N__23491\
        );

    \I__5108\ : LocalMux
    port map (
            O => \N__23491\,
            I => \N__23488\
        );

    \I__5107\ : Span4Mux_s2_h
    port map (
            O => \N__23488\,
            I => \N__23485\
        );

    \I__5106\ : Odrv4
    port map (
            O => \N__23485\,
            I => led_c_2
        );

    \I__5105\ : InMux
    port map (
            O => \N__23482\,
            I => \N__23479\
        );

    \I__5104\ : LocalMux
    port map (
            O => \N__23479\,
            I => \N__23473\
        );

    \I__5103\ : InMux
    port map (
            O => \N__23478\,
            I => \N__23470\
        );

    \I__5102\ : InMux
    port map (
            O => \N__23477\,
            I => \N__23465\
        );

    \I__5101\ : InMux
    port map (
            O => \N__23476\,
            I => \N__23465\
        );

    \I__5100\ : Odrv4
    port map (
            O => \N__23473\,
            I => \Lab_UT.dictrl.r_Sone_init5\
        );

    \I__5099\ : LocalMux
    port map (
            O => \N__23470\,
            I => \Lab_UT.dictrl.r_Sone_init5\
        );

    \I__5098\ : LocalMux
    port map (
            O => \N__23465\,
            I => \Lab_UT.dictrl.r_Sone_init5\
        );

    \I__5097\ : CascadeMux
    port map (
            O => \N__23458\,
            I => \N__23449\
        );

    \I__5096\ : CascadeMux
    port map (
            O => \N__23457\,
            I => \N__23441\
        );

    \I__5095\ : InMux
    port map (
            O => \N__23456\,
            I => \N__23432\
        );

    \I__5094\ : InMux
    port map (
            O => \N__23455\,
            I => \N__23423\
        );

    \I__5093\ : InMux
    port map (
            O => \N__23454\,
            I => \N__23423\
        );

    \I__5092\ : InMux
    port map (
            O => \N__23453\,
            I => \N__23423\
        );

    \I__5091\ : InMux
    port map (
            O => \N__23452\,
            I => \N__23415\
        );

    \I__5090\ : InMux
    port map (
            O => \N__23449\,
            I => \N__23415\
        );

    \I__5089\ : InMux
    port map (
            O => \N__23448\,
            I => \N__23415\
        );

    \I__5088\ : InMux
    port map (
            O => \N__23447\,
            I => \N__23412\
        );

    \I__5087\ : InMux
    port map (
            O => \N__23446\,
            I => \N__23405\
        );

    \I__5086\ : InMux
    port map (
            O => \N__23445\,
            I => \N__23405\
        );

    \I__5085\ : InMux
    port map (
            O => \N__23444\,
            I => \N__23405\
        );

    \I__5084\ : InMux
    port map (
            O => \N__23441\,
            I => \N__23402\
        );

    \I__5083\ : InMux
    port map (
            O => \N__23440\,
            I => \N__23397\
        );

    \I__5082\ : InMux
    port map (
            O => \N__23439\,
            I => \N__23397\
        );

    \I__5081\ : InMux
    port map (
            O => \N__23438\,
            I => \N__23390\
        );

    \I__5080\ : InMux
    port map (
            O => \N__23437\,
            I => \N__23390\
        );

    \I__5079\ : InMux
    port map (
            O => \N__23436\,
            I => \N__23390\
        );

    \I__5078\ : InMux
    port map (
            O => \N__23435\,
            I => \N__23385\
        );

    \I__5077\ : LocalMux
    port map (
            O => \N__23432\,
            I => \N__23382\
        );

    \I__5076\ : InMux
    port map (
            O => \N__23431\,
            I => \N__23378\
        );

    \I__5075\ : InMux
    port map (
            O => \N__23430\,
            I => \N__23372\
        );

    \I__5074\ : LocalMux
    port map (
            O => \N__23423\,
            I => \N__23369\
        );

    \I__5073\ : InMux
    port map (
            O => \N__23422\,
            I => \N__23366\
        );

    \I__5072\ : LocalMux
    port map (
            O => \N__23415\,
            I => \N__23363\
        );

    \I__5071\ : LocalMux
    port map (
            O => \N__23412\,
            I => \N__23358\
        );

    \I__5070\ : LocalMux
    port map (
            O => \N__23405\,
            I => \N__23358\
        );

    \I__5069\ : LocalMux
    port map (
            O => \N__23402\,
            I => \N__23351\
        );

    \I__5068\ : LocalMux
    port map (
            O => \N__23397\,
            I => \N__23351\
        );

    \I__5067\ : LocalMux
    port map (
            O => \N__23390\,
            I => \N__23351\
        );

    \I__5066\ : InMux
    port map (
            O => \N__23389\,
            I => \N__23346\
        );

    \I__5065\ : InMux
    port map (
            O => \N__23388\,
            I => \N__23346\
        );

    \I__5064\ : LocalMux
    port map (
            O => \N__23385\,
            I => \N__23337\
        );

    \I__5063\ : Span4Mux_s3_h
    port map (
            O => \N__23382\,
            I => \N__23334\
        );

    \I__5062\ : InMux
    port map (
            O => \N__23381\,
            I => \N__23331\
        );

    \I__5061\ : LocalMux
    port map (
            O => \N__23378\,
            I => \N__23328\
        );

    \I__5060\ : InMux
    port map (
            O => \N__23377\,
            I => \N__23321\
        );

    \I__5059\ : InMux
    port map (
            O => \N__23376\,
            I => \N__23321\
        );

    \I__5058\ : InMux
    port map (
            O => \N__23375\,
            I => \N__23318\
        );

    \I__5057\ : LocalMux
    port map (
            O => \N__23372\,
            I => \N__23315\
        );

    \I__5056\ : Span4Mux_v
    port map (
            O => \N__23369\,
            I => \N__23308\
        );

    \I__5055\ : LocalMux
    port map (
            O => \N__23366\,
            I => \N__23308\
        );

    \I__5054\ : Span4Mux_h
    port map (
            O => \N__23363\,
            I => \N__23308\
        );

    \I__5053\ : Span4Mux_v
    port map (
            O => \N__23358\,
            I => \N__23301\
        );

    \I__5052\ : Span4Mux_h
    port map (
            O => \N__23351\,
            I => \N__23301\
        );

    \I__5051\ : LocalMux
    port map (
            O => \N__23346\,
            I => \N__23301\
        );

    \I__5050\ : InMux
    port map (
            O => \N__23345\,
            I => \N__23298\
        );

    \I__5049\ : InMux
    port map (
            O => \N__23344\,
            I => \N__23295\
        );

    \I__5048\ : InMux
    port map (
            O => \N__23343\,
            I => \N__23286\
        );

    \I__5047\ : InMux
    port map (
            O => \N__23342\,
            I => \N__23286\
        );

    \I__5046\ : InMux
    port map (
            O => \N__23341\,
            I => \N__23286\
        );

    \I__5045\ : InMux
    port map (
            O => \N__23340\,
            I => \N__23286\
        );

    \I__5044\ : Span4Mux_h
    port map (
            O => \N__23337\,
            I => \N__23277\
        );

    \I__5043\ : Span4Mux_h
    port map (
            O => \N__23334\,
            I => \N__23277\
        );

    \I__5042\ : LocalMux
    port map (
            O => \N__23331\,
            I => \N__23277\
        );

    \I__5041\ : Span4Mux_v
    port map (
            O => \N__23328\,
            I => \N__23277\
        );

    \I__5040\ : InMux
    port map (
            O => \N__23327\,
            I => \N__23272\
        );

    \I__5039\ : InMux
    port map (
            O => \N__23326\,
            I => \N__23272\
        );

    \I__5038\ : LocalMux
    port map (
            O => \N__23321\,
            I => \N__23261\
        );

    \I__5037\ : LocalMux
    port map (
            O => \N__23318\,
            I => \N__23261\
        );

    \I__5036\ : Span4Mux_h
    port map (
            O => \N__23315\,
            I => \N__23261\
        );

    \I__5035\ : Span4Mux_h
    port map (
            O => \N__23308\,
            I => \N__23261\
        );

    \I__5034\ : Span4Mux_h
    port map (
            O => \N__23301\,
            I => \N__23261\
        );

    \I__5033\ : LocalMux
    port map (
            O => \N__23298\,
            I => \Lab_UT_dictrl_r_Sone_init17\
        );

    \I__5032\ : LocalMux
    port map (
            O => \N__23295\,
            I => \Lab_UT_dictrl_r_Sone_init17\
        );

    \I__5031\ : LocalMux
    port map (
            O => \N__23286\,
            I => \Lab_UT_dictrl_r_Sone_init17\
        );

    \I__5030\ : Odrv4
    port map (
            O => \N__23277\,
            I => \Lab_UT_dictrl_r_Sone_init17\
        );

    \I__5029\ : LocalMux
    port map (
            O => \N__23272\,
            I => \Lab_UT_dictrl_r_Sone_init17\
        );

    \I__5028\ : Odrv4
    port map (
            O => \N__23261\,
            I => \Lab_UT_dictrl_r_Sone_init17\
        );

    \I__5027\ : InMux
    port map (
            O => \N__23248\,
            I => \N__23241\
        );

    \I__5026\ : InMux
    port map (
            O => \N__23247\,
            I => \N__23241\
        );

    \I__5025\ : InMux
    port map (
            O => \N__23246\,
            I => \N__23236\
        );

    \I__5024\ : LocalMux
    port map (
            O => \N__23241\,
            I => \N__23229\
        );

    \I__5023\ : InMux
    port map (
            O => \N__23240\,
            I => \N__23224\
        );

    \I__5022\ : InMux
    port map (
            O => \N__23239\,
            I => \N__23224\
        );

    \I__5021\ : LocalMux
    port map (
            O => \N__23236\,
            I => \N__23217\
        );

    \I__5020\ : InMux
    port map (
            O => \N__23235\,
            I => \N__23214\
        );

    \I__5019\ : InMux
    port map (
            O => \N__23234\,
            I => \N__23207\
        );

    \I__5018\ : InMux
    port map (
            O => \N__23233\,
            I => \N__23207\
        );

    \I__5017\ : InMux
    port map (
            O => \N__23232\,
            I => \N__23207\
        );

    \I__5016\ : Span4Mux_s1_v
    port map (
            O => \N__23229\,
            I => \N__23202\
        );

    \I__5015\ : LocalMux
    port map (
            O => \N__23224\,
            I => \N__23202\
        );

    \I__5014\ : InMux
    port map (
            O => \N__23223\,
            I => \N__23199\
        );

    \I__5013\ : InMux
    port map (
            O => \N__23222\,
            I => \N__23192\
        );

    \I__5012\ : InMux
    port map (
            O => \N__23221\,
            I => \N__23192\
        );

    \I__5011\ : InMux
    port map (
            O => \N__23220\,
            I => \N__23192\
        );

    \I__5010\ : Span4Mux_v
    port map (
            O => \N__23217\,
            I => \N__23187\
        );

    \I__5009\ : LocalMux
    port map (
            O => \N__23214\,
            I => \N__23187\
        );

    \I__5008\ : LocalMux
    port map (
            O => \N__23207\,
            I => \Lab_UT.uu0.un4_l_count_0\
        );

    \I__5007\ : Odrv4
    port map (
            O => \N__23202\,
            I => \Lab_UT.uu0.un4_l_count_0\
        );

    \I__5006\ : LocalMux
    port map (
            O => \N__23199\,
            I => \Lab_UT.uu0.un4_l_count_0\
        );

    \I__5005\ : LocalMux
    port map (
            O => \N__23192\,
            I => \Lab_UT.uu0.un4_l_count_0\
        );

    \I__5004\ : Odrv4
    port map (
            O => \N__23187\,
            I => \Lab_UT.uu0.un4_l_count_0\
        );

    \I__5003\ : CascadeMux
    port map (
            O => \N__23176\,
            I => \N__23171\
        );

    \I__5002\ : InMux
    port map (
            O => \N__23175\,
            I => \N__23163\
        );

    \I__5001\ : InMux
    port map (
            O => \N__23174\,
            I => \N__23163\
        );

    \I__5000\ : InMux
    port map (
            O => \N__23171\,
            I => \N__23163\
        );

    \I__4999\ : CascadeMux
    port map (
            O => \N__23170\,
            I => \N__23158\
        );

    \I__4998\ : LocalMux
    port map (
            O => \N__23163\,
            I => \N__23154\
        );

    \I__4997\ : InMux
    port map (
            O => \N__23162\,
            I => \N__23147\
        );

    \I__4996\ : InMux
    port map (
            O => \N__23161\,
            I => \N__23147\
        );

    \I__4995\ : InMux
    port map (
            O => \N__23158\,
            I => \N__23147\
        );

    \I__4994\ : InMux
    port map (
            O => \N__23157\,
            I => \N__23144\
        );

    \I__4993\ : Span4Mux_h
    port map (
            O => \N__23154\,
            I => \N__23141\
        );

    \I__4992\ : LocalMux
    port map (
            O => \N__23147\,
            I => \N__23138\
        );

    \I__4991\ : LocalMux
    port map (
            O => \N__23144\,
            I => \Lab_UT.halfPulse\
        );

    \I__4990\ : Odrv4
    port map (
            O => \N__23141\,
            I => \Lab_UT.halfPulse\
        );

    \I__4989\ : Odrv4
    port map (
            O => \N__23138\,
            I => \Lab_UT.halfPulse\
        );

    \I__4988\ : InMux
    port map (
            O => \N__23131\,
            I => \N__23127\
        );

    \I__4987\ : InMux
    port map (
            O => \N__23130\,
            I => \N__23124\
        );

    \I__4986\ : LocalMux
    port map (
            O => \N__23127\,
            I => \N__23121\
        );

    \I__4985\ : LocalMux
    port map (
            O => \N__23124\,
            I => \N__23118\
        );

    \I__4984\ : Odrv12
    port map (
            O => \N__23121\,
            I => \Lab_UT.displayAlarmZ0Z_1\
        );

    \I__4983\ : Odrv4
    port map (
            O => \N__23118\,
            I => \Lab_UT.displayAlarmZ0Z_1\
        );

    \I__4982\ : CascadeMux
    port map (
            O => \N__23113\,
            I => \N__23109\
        );

    \I__4981\ : CascadeMux
    port map (
            O => \N__23112\,
            I => \N__23106\
        );

    \I__4980\ : InMux
    port map (
            O => \N__23109\,
            I => \N__23102\
        );

    \I__4979\ : InMux
    port map (
            O => \N__23106\,
            I => \N__23097\
        );

    \I__4978\ : InMux
    port map (
            O => \N__23105\,
            I => \N__23097\
        );

    \I__4977\ : LocalMux
    port map (
            O => \N__23102\,
            I => \Lab_UT.dicLdStens\
        );

    \I__4976\ : LocalMux
    port map (
            O => \N__23097\,
            I => \Lab_UT.dicLdStens\
        );

    \I__4975\ : InMux
    port map (
            O => \N__23092\,
            I => \N__23087\
        );

    \I__4974\ : InMux
    port map (
            O => \N__23091\,
            I => \N__23082\
        );

    \I__4973\ : InMux
    port map (
            O => \N__23090\,
            I => \N__23082\
        );

    \I__4972\ : LocalMux
    port map (
            O => \N__23087\,
            I => \Lab_UT.dicLdStens_latmux\
        );

    \I__4971\ : LocalMux
    port map (
            O => \N__23082\,
            I => \Lab_UT.dicLdStens_latmux\
        );

    \I__4970\ : InMux
    port map (
            O => \N__23077\,
            I => \N__23072\
        );

    \I__4969\ : InMux
    port map (
            O => \N__23076\,
            I => \N__23069\
        );

    \I__4968\ : InMux
    port map (
            O => \N__23075\,
            I => \N__23066\
        );

    \I__4967\ : LocalMux
    port map (
            O => \N__23072\,
            I => \Lab_UT.di_ASones_0\
        );

    \I__4966\ : LocalMux
    port map (
            O => \N__23069\,
            I => \Lab_UT.di_ASones_0\
        );

    \I__4965\ : LocalMux
    port map (
            O => \N__23066\,
            I => \Lab_UT.di_ASones_0\
        );

    \I__4964\ : InMux
    port map (
            O => \N__23059\,
            I => \N__23054\
        );

    \I__4963\ : InMux
    port map (
            O => \N__23058\,
            I => \N__23051\
        );

    \I__4962\ : InMux
    port map (
            O => \N__23057\,
            I => \N__23048\
        );

    \I__4961\ : LocalMux
    port map (
            O => \N__23054\,
            I => \N__23045\
        );

    \I__4960\ : LocalMux
    port map (
            O => \N__23051\,
            I => \Lab_UT.di_ASones_1\
        );

    \I__4959\ : LocalMux
    port map (
            O => \N__23048\,
            I => \Lab_UT.di_ASones_1\
        );

    \I__4958\ : Odrv4
    port map (
            O => \N__23045\,
            I => \Lab_UT.di_ASones_1\
        );

    \I__4957\ : InMux
    port map (
            O => \N__23038\,
            I => \N__23033\
        );

    \I__4956\ : InMux
    port map (
            O => \N__23037\,
            I => \N__23030\
        );

    \I__4955\ : InMux
    port map (
            O => \N__23036\,
            I => \N__23027\
        );

    \I__4954\ : LocalMux
    port map (
            O => \N__23033\,
            I => \Lab_UT.di_ASones_2\
        );

    \I__4953\ : LocalMux
    port map (
            O => \N__23030\,
            I => \Lab_UT.di_ASones_2\
        );

    \I__4952\ : LocalMux
    port map (
            O => \N__23027\,
            I => \Lab_UT.di_ASones_2\
        );

    \I__4951\ : CascadeMux
    port map (
            O => \N__23020\,
            I => \N__23015\
        );

    \I__4950\ : InMux
    port map (
            O => \N__23019\,
            I => \N__23011\
        );

    \I__4949\ : InMux
    port map (
            O => \N__23018\,
            I => \N__23008\
        );

    \I__4948\ : InMux
    port map (
            O => \N__23015\,
            I => \N__23003\
        );

    \I__4947\ : InMux
    port map (
            O => \N__23014\,
            I => \N__23003\
        );

    \I__4946\ : LocalMux
    port map (
            O => \N__23011\,
            I => \N__22998\
        );

    \I__4945\ : LocalMux
    port map (
            O => \N__23008\,
            I => \N__22998\
        );

    \I__4944\ : LocalMux
    port map (
            O => \N__23003\,
            I => \N__22995\
        );

    \I__4943\ : Span4Mux_h
    port map (
            O => \N__22998\,
            I => \N__22992\
        );

    \I__4942\ : Span4Mux_h
    port map (
            O => \N__22995\,
            I => \N__22989\
        );

    \I__4941\ : Odrv4
    port map (
            O => \N__22992\,
            I => \Lab_UT.ld_enable_AMtens\
        );

    \I__4940\ : Odrv4
    port map (
            O => \N__22989\,
            I => \Lab_UT.ld_enable_AMtens\
        );

    \I__4939\ : InMux
    port map (
            O => \N__22984\,
            I => \N__22980\
        );

    \I__4938\ : InMux
    port map (
            O => \N__22983\,
            I => \N__22976\
        );

    \I__4937\ : LocalMux
    port map (
            O => \N__22980\,
            I => \N__22973\
        );

    \I__4936\ : InMux
    port map (
            O => \N__22979\,
            I => \N__22970\
        );

    \I__4935\ : LocalMux
    port map (
            O => \N__22976\,
            I => \Lab_UT.di_AStens_3\
        );

    \I__4934\ : Odrv4
    port map (
            O => \N__22973\,
            I => \Lab_UT.di_AStens_3\
        );

    \I__4933\ : LocalMux
    port map (
            O => \N__22970\,
            I => \Lab_UT.di_AStens_3\
        );

    \I__4932\ : InMux
    port map (
            O => \N__22963\,
            I => \N__22954\
        );

    \I__4931\ : InMux
    port map (
            O => \N__22962\,
            I => \N__22954\
        );

    \I__4930\ : InMux
    port map (
            O => \N__22961\,
            I => \N__22954\
        );

    \I__4929\ : LocalMux
    port map (
            O => \N__22954\,
            I => \N__22950\
        );

    \I__4928\ : InMux
    port map (
            O => \N__22953\,
            I => \N__22947\
        );

    \I__4927\ : Span4Mux_v
    port map (
            O => \N__22950\,
            I => \N__22944\
        );

    \I__4926\ : LocalMux
    port map (
            O => \N__22947\,
            I => \N__22941\
        );

    \I__4925\ : Span4Mux_v
    port map (
            O => \N__22944\,
            I => \N__22938\
        );

    \I__4924\ : Span4Mux_h
    port map (
            O => \N__22941\,
            I => \N__22935\
        );

    \I__4923\ : Odrv4
    port map (
            O => \N__22938\,
            I => \Lab_UT.ld_enable_ASones\
        );

    \I__4922\ : Odrv4
    port map (
            O => \N__22935\,
            I => \Lab_UT.ld_enable_ASones\
        );

    \I__4921\ : InMux
    port map (
            O => \N__22930\,
            I => \N__22926\
        );

    \I__4920\ : InMux
    port map (
            O => \N__22929\,
            I => \N__22922\
        );

    \I__4919\ : LocalMux
    port map (
            O => \N__22926\,
            I => \N__22919\
        );

    \I__4918\ : InMux
    port map (
            O => \N__22925\,
            I => \N__22916\
        );

    \I__4917\ : LocalMux
    port map (
            O => \N__22922\,
            I => \Lab_UT.di_ASones_3\
        );

    \I__4916\ : Odrv4
    port map (
            O => \N__22919\,
            I => \Lab_UT.di_ASones_3\
        );

    \I__4915\ : LocalMux
    port map (
            O => \N__22916\,
            I => \Lab_UT.di_ASones_3\
        );

    \I__4914\ : InMux
    port map (
            O => \N__22909\,
            I => \N__22897\
        );

    \I__4913\ : InMux
    port map (
            O => \N__22908\,
            I => \N__22897\
        );

    \I__4912\ : InMux
    port map (
            O => \N__22907\,
            I => \N__22897\
        );

    \I__4911\ : InMux
    port map (
            O => \N__22906\,
            I => \N__22897\
        );

    \I__4910\ : LocalMux
    port map (
            O => \N__22897\,
            I => \N__22894\
        );

    \I__4909\ : Span4Mux_v
    port map (
            O => \N__22894\,
            I => \N__22891\
        );

    \I__4908\ : Odrv4
    port map (
            O => \N__22891\,
            I => \Lab_UT.ld_enable_AStens\
        );

    \I__4907\ : InMux
    port map (
            O => \N__22888\,
            I => \N__22885\
        );

    \I__4906\ : LocalMux
    port map (
            O => \N__22885\,
            I => \Lab_UT.display.dOutP_0_iv_i_1_1\
        );

    \I__4905\ : CascadeMux
    port map (
            O => \N__22882\,
            I => \N__22878\
        );

    \I__4904\ : CascadeMux
    port map (
            O => \N__22881\,
            I => \N__22875\
        );

    \I__4903\ : InMux
    port map (
            O => \N__22878\,
            I => \N__22864\
        );

    \I__4902\ : InMux
    port map (
            O => \N__22875\,
            I => \N__22864\
        );

    \I__4901\ : InMux
    port map (
            O => \N__22874\,
            I => \N__22864\
        );

    \I__4900\ : InMux
    port map (
            O => \N__22873\,
            I => \N__22864\
        );

    \I__4899\ : LocalMux
    port map (
            O => \N__22864\,
            I => \Lab_UT.display.N_150\
        );

    \I__4898\ : CascadeMux
    port map (
            O => \N__22861\,
            I => \Lab_UT.display.N_101_cascade_\
        );

    \I__4897\ : InMux
    port map (
            O => \N__22858\,
            I => \N__22855\
        );

    \I__4896\ : LocalMux
    port map (
            O => \N__22855\,
            I => \N__22851\
        );

    \I__4895\ : InMux
    port map (
            O => \N__22854\,
            I => \N__22848\
        );

    \I__4894\ : Odrv4
    port map (
            O => \N__22851\,
            I => \Lab_UT.display.N_88\
        );

    \I__4893\ : LocalMux
    port map (
            O => \N__22848\,
            I => \Lab_UT.display.N_88\
        );

    \I__4892\ : CascadeMux
    port map (
            O => \N__22843\,
            I => \Lab_UT.display.dOutP_0_iv_i_0_3_cascade_\
        );

    \I__4891\ : InMux
    port map (
            O => \N__22840\,
            I => \N__22837\
        );

    \I__4890\ : LocalMux
    port map (
            O => \N__22837\,
            I => \Lab_UT.display.dOutP_0_iv_i_2_3\
        );

    \I__4889\ : InMux
    port map (
            O => \N__22834\,
            I => \N__22831\
        );

    \I__4888\ : LocalMux
    port map (
            O => \N__22831\,
            I => \N__22828\
        );

    \I__4887\ : Span4Mux_v
    port map (
            O => \N__22828\,
            I => \N__22824\
        );

    \I__4886\ : InMux
    port map (
            O => \N__22827\,
            I => \N__22821\
        );

    \I__4885\ : Span4Mux_h
    port map (
            O => \N__22824\,
            I => \N__22815\
        );

    \I__4884\ : LocalMux
    port map (
            O => \N__22821\,
            I => \N__22815\
        );

    \I__4883\ : InMux
    port map (
            O => \N__22820\,
            I => \N__22812\
        );

    \I__4882\ : Odrv4
    port map (
            O => \N__22815\,
            I => \L3_tx_data_3\
        );

    \I__4881\ : LocalMux
    port map (
            O => \N__22812\,
            I => \L3_tx_data_3\
        );

    \I__4880\ : InMux
    port map (
            O => \N__22807\,
            I => \N__22803\
        );

    \I__4879\ : CascadeMux
    port map (
            O => \N__22806\,
            I => \N__22800\
        );

    \I__4878\ : LocalMux
    port map (
            O => \N__22803\,
            I => \N__22797\
        );

    \I__4877\ : InMux
    port map (
            O => \N__22800\,
            I => \N__22794\
        );

    \I__4876\ : Span4Mux_h
    port map (
            O => \N__22797\,
            I => \N__22787\
        );

    \I__4875\ : LocalMux
    port map (
            O => \N__22794\,
            I => \N__22787\
        );

    \I__4874\ : InMux
    port map (
            O => \N__22793\,
            I => \N__22784\
        );

    \I__4873\ : CascadeMux
    port map (
            O => \N__22792\,
            I => \N__22781\
        );

    \I__4872\ : Span4Mux_h
    port map (
            O => \N__22787\,
            I => \N__22776\
        );

    \I__4871\ : LocalMux
    port map (
            O => \N__22784\,
            I => \N__22776\
        );

    \I__4870\ : InMux
    port map (
            O => \N__22781\,
            I => \N__22773\
        );

    \I__4869\ : Span4Mux_h
    port map (
            O => \N__22776\,
            I => \N__22770\
        );

    \I__4868\ : LocalMux
    port map (
            O => \N__22773\,
            I => \uu2.r_addrZ0Z_5\
        );

    \I__4867\ : Odrv4
    port map (
            O => \N__22770\,
            I => \uu2.r_addrZ0Z_5\
        );

    \I__4866\ : InMux
    port map (
            O => \N__22765\,
            I => \N__22761\
        );

    \I__4865\ : CascadeMux
    port map (
            O => \N__22764\,
            I => \N__22757\
        );

    \I__4864\ : LocalMux
    port map (
            O => \N__22761\,
            I => \N__22754\
        );

    \I__4863\ : InMux
    port map (
            O => \N__22760\,
            I => \N__22751\
        );

    \I__4862\ : InMux
    port map (
            O => \N__22757\,
            I => \N__22748\
        );

    \I__4861\ : Span4Mux_h
    port map (
            O => \N__22754\,
            I => \N__22745\
        );

    \I__4860\ : LocalMux
    port map (
            O => \N__22751\,
            I => \Lab_UT.di_AMones_0\
        );

    \I__4859\ : LocalMux
    port map (
            O => \N__22748\,
            I => \Lab_UT.di_AMones_0\
        );

    \I__4858\ : Odrv4
    port map (
            O => \N__22745\,
            I => \Lab_UT.di_AMones_0\
        );

    \I__4857\ : InMux
    port map (
            O => \N__22738\,
            I => \N__22735\
        );

    \I__4856\ : LocalMux
    port map (
            O => \N__22735\,
            I => \N__22730\
        );

    \I__4855\ : InMux
    port map (
            O => \N__22734\,
            I => \N__22727\
        );

    \I__4854\ : InMux
    port map (
            O => \N__22733\,
            I => \N__22724\
        );

    \I__4853\ : Span4Mux_v
    port map (
            O => \N__22730\,
            I => \N__22721\
        );

    \I__4852\ : LocalMux
    port map (
            O => \N__22727\,
            I => \Lab_UT.di_AMones_2\
        );

    \I__4851\ : LocalMux
    port map (
            O => \N__22724\,
            I => \Lab_UT.di_AMones_2\
        );

    \I__4850\ : Odrv4
    port map (
            O => \N__22721\,
            I => \Lab_UT.di_AMones_2\
        );

    \I__4849\ : InMux
    port map (
            O => \N__22714\,
            I => \N__22702\
        );

    \I__4848\ : InMux
    port map (
            O => \N__22713\,
            I => \N__22702\
        );

    \I__4847\ : InMux
    port map (
            O => \N__22712\,
            I => \N__22702\
        );

    \I__4846\ : InMux
    port map (
            O => \N__22711\,
            I => \N__22702\
        );

    \I__4845\ : LocalMux
    port map (
            O => \N__22702\,
            I => \N__22699\
        );

    \I__4844\ : Span4Mux_v
    port map (
            O => \N__22699\,
            I => \N__22696\
        );

    \I__4843\ : Odrv4
    port map (
            O => \N__22696\,
            I => \Lab_UT.ld_enable_AMones\
        );

    \I__4842\ : InMux
    port map (
            O => \N__22693\,
            I => \N__22690\
        );

    \I__4841\ : LocalMux
    port map (
            O => \N__22690\,
            I => \N__22685\
        );

    \I__4840\ : InMux
    port map (
            O => \N__22689\,
            I => \N__22682\
        );

    \I__4839\ : InMux
    port map (
            O => \N__22688\,
            I => \N__22679\
        );

    \I__4838\ : Span4Mux_h
    port map (
            O => \N__22685\,
            I => \N__22676\
        );

    \I__4837\ : LocalMux
    port map (
            O => \N__22682\,
            I => \Lab_UT.di_AMones_3\
        );

    \I__4836\ : LocalMux
    port map (
            O => \N__22679\,
            I => \Lab_UT.di_AMones_3\
        );

    \I__4835\ : Odrv4
    port map (
            O => \N__22676\,
            I => \Lab_UT.di_AMones_3\
        );

    \I__4834\ : CascadeMux
    port map (
            O => \N__22669\,
            I => \Lab_UT.display.N_88_cascade_\
        );

    \I__4833\ : InMux
    port map (
            O => \N__22666\,
            I => \N__22662\
        );

    \I__4832\ : CascadeMux
    port map (
            O => \N__22665\,
            I => \N__22658\
        );

    \I__4831\ : LocalMux
    port map (
            O => \N__22662\,
            I => \N__22655\
        );

    \I__4830\ : InMux
    port map (
            O => \N__22661\,
            I => \N__22652\
        );

    \I__4829\ : InMux
    port map (
            O => \N__22658\,
            I => \N__22649\
        );

    \I__4828\ : Odrv12
    port map (
            O => \N__22655\,
            I => \L3_tx_data_1\
        );

    \I__4827\ : LocalMux
    port map (
            O => \N__22652\,
            I => \L3_tx_data_1\
        );

    \I__4826\ : LocalMux
    port map (
            O => \N__22649\,
            I => \L3_tx_data_1\
        );

    \I__4825\ : CascadeMux
    port map (
            O => \N__22642\,
            I => \Lab_UT.display.N_120_cascade_\
        );

    \I__4824\ : InMux
    port map (
            O => \N__22639\,
            I => \N__22636\
        );

    \I__4823\ : LocalMux
    port map (
            O => \N__22636\,
            I => \N__22633\
        );

    \I__4822\ : Span4Mux_h
    port map (
            O => \N__22633\,
            I => \N__22628\
        );

    \I__4821\ : InMux
    port map (
            O => \N__22632\,
            I => \N__22623\
        );

    \I__4820\ : InMux
    port map (
            O => \N__22631\,
            I => \N__22623\
        );

    \I__4819\ : Odrv4
    port map (
            O => \N__22628\,
            I => \L3_tx_data_4\
        );

    \I__4818\ : LocalMux
    port map (
            O => \N__22623\,
            I => \L3_tx_data_4\
        );

    \I__4817\ : InMux
    port map (
            O => \N__22618\,
            I => \N__22615\
        );

    \I__4816\ : LocalMux
    port map (
            O => \N__22615\,
            I => \N__22610\
        );

    \I__4815\ : InMux
    port map (
            O => \N__22614\,
            I => \N__22605\
        );

    \I__4814\ : InMux
    port map (
            O => \N__22613\,
            I => \N__22605\
        );

    \I__4813\ : Odrv12
    port map (
            O => \N__22610\,
            I => \L3_tx_data_5\
        );

    \I__4812\ : LocalMux
    port map (
            O => \N__22605\,
            I => \L3_tx_data_5\
        );

    \I__4811\ : CascadeMux
    port map (
            O => \N__22600\,
            I => \Lab_UT.display.N_153_cascade_\
        );

    \I__4810\ : InMux
    port map (
            O => \N__22597\,
            I => \N__22582\
        );

    \I__4809\ : InMux
    port map (
            O => \N__22596\,
            I => \N__22582\
        );

    \I__4808\ : InMux
    port map (
            O => \N__22595\,
            I => \N__22582\
        );

    \I__4807\ : InMux
    port map (
            O => \N__22594\,
            I => \N__22582\
        );

    \I__4806\ : InMux
    port map (
            O => \N__22593\,
            I => \N__22582\
        );

    \I__4805\ : LocalMux
    port map (
            O => \N__22582\,
            I => \Lab_UT.uu0.l_precountZ0Z_1\
        );

    \I__4804\ : InMux
    port map (
            O => \N__22579\,
            I => \N__22569\
        );

    \I__4803\ : InMux
    port map (
            O => \N__22578\,
            I => \N__22569\
        );

    \I__4802\ : InMux
    port map (
            O => \N__22577\,
            I => \N__22569\
        );

    \I__4801\ : InMux
    port map (
            O => \N__22576\,
            I => \N__22566\
        );

    \I__4800\ : LocalMux
    port map (
            O => \N__22569\,
            I => \Lab_UT.uu0.l_countZ0Z_16\
        );

    \I__4799\ : LocalMux
    port map (
            O => \N__22566\,
            I => \Lab_UT.uu0.l_countZ0Z_16\
        );

    \I__4798\ : CascadeMux
    port map (
            O => \N__22561\,
            I => \N__22557\
        );

    \I__4797\ : InMux
    port map (
            O => \N__22560\,
            I => \N__22551\
        );

    \I__4796\ : InMux
    port map (
            O => \N__22557\,
            I => \N__22551\
        );

    \I__4795\ : InMux
    port map (
            O => \N__22556\,
            I => \N__22548\
        );

    \I__4794\ : LocalMux
    port map (
            O => \N__22551\,
            I => \N__22543\
        );

    \I__4793\ : LocalMux
    port map (
            O => \N__22548\,
            I => \N__22543\
        );

    \I__4792\ : Odrv4
    port map (
            O => \N__22543\,
            I => \Lab_UT.uu0.l_countZ0Z_11\
        );

    \I__4791\ : CascadeMux
    port map (
            O => \N__22540\,
            I => \N__22534\
        );

    \I__4790\ : InMux
    port map (
            O => \N__22539\,
            I => \N__22525\
        );

    \I__4789\ : InMux
    port map (
            O => \N__22538\,
            I => \N__22525\
        );

    \I__4788\ : InMux
    port map (
            O => \N__22537\,
            I => \N__22525\
        );

    \I__4787\ : InMux
    port map (
            O => \N__22534\,
            I => \N__22525\
        );

    \I__4786\ : LocalMux
    port map (
            O => \N__22525\,
            I => \Lab_UT.uu0.l_precountZ0Z_2\
        );

    \I__4785\ : CascadeMux
    port map (
            O => \N__22522\,
            I => \N__22516\
        );

    \I__4784\ : InMux
    port map (
            O => \N__22521\,
            I => \N__22506\
        );

    \I__4783\ : InMux
    port map (
            O => \N__22520\,
            I => \N__22506\
        );

    \I__4782\ : InMux
    port map (
            O => \N__22519\,
            I => \N__22506\
        );

    \I__4781\ : InMux
    port map (
            O => \N__22516\,
            I => \N__22506\
        );

    \I__4780\ : InMux
    port map (
            O => \N__22515\,
            I => \N__22503\
        );

    \I__4779\ : LocalMux
    port map (
            O => \N__22506\,
            I => \Lab_UT.uu0.l_countZ0Z_0\
        );

    \I__4778\ : LocalMux
    port map (
            O => \N__22503\,
            I => \Lab_UT.uu0.l_countZ0Z_0\
        );

    \I__4777\ : InMux
    port map (
            O => \N__22498\,
            I => \N__22495\
        );

    \I__4776\ : LocalMux
    port map (
            O => \N__22495\,
            I => \Lab_UT.uu0.un4_l_count_13\
        );

    \I__4775\ : CascadeMux
    port map (
            O => \N__22492\,
            I => \N__22489\
        );

    \I__4774\ : InMux
    port map (
            O => \N__22489\,
            I => \N__22481\
        );

    \I__4773\ : InMux
    port map (
            O => \N__22488\,
            I => \N__22481\
        );

    \I__4772\ : InMux
    port map (
            O => \N__22487\,
            I => \N__22478\
        );

    \I__4771\ : InMux
    port map (
            O => \N__22486\,
            I => \N__22475\
        );

    \I__4770\ : LocalMux
    port map (
            O => \N__22481\,
            I => \N__22472\
        );

    \I__4769\ : LocalMux
    port map (
            O => \N__22478\,
            I => \N__22469\
        );

    \I__4768\ : LocalMux
    port map (
            O => \N__22475\,
            I => \uu2.w_addr_userZ0Z_5\
        );

    \I__4767\ : Odrv12
    port map (
            O => \N__22472\,
            I => \uu2.w_addr_userZ0Z_5\
        );

    \I__4766\ : Odrv4
    port map (
            O => \N__22469\,
            I => \uu2.w_addr_userZ0Z_5\
        );

    \I__4765\ : CascadeMux
    port map (
            O => \N__22462\,
            I => \N__22456\
        );

    \I__4764\ : InMux
    port map (
            O => \N__22461\,
            I => \N__22450\
        );

    \I__4763\ : InMux
    port map (
            O => \N__22460\,
            I => \N__22450\
        );

    \I__4762\ : InMux
    port map (
            O => \N__22459\,
            I => \N__22447\
        );

    \I__4761\ : InMux
    port map (
            O => \N__22456\,
            I => \N__22442\
        );

    \I__4760\ : InMux
    port map (
            O => \N__22455\,
            I => \N__22442\
        );

    \I__4759\ : LocalMux
    port map (
            O => \N__22450\,
            I => \N__22439\
        );

    \I__4758\ : LocalMux
    port map (
            O => \N__22447\,
            I => \N__22436\
        );

    \I__4757\ : LocalMux
    port map (
            O => \N__22442\,
            I => \uu2.w_addr_userZ0Z_4\
        );

    \I__4756\ : Odrv12
    port map (
            O => \N__22439\,
            I => \uu2.w_addr_userZ0Z_4\
        );

    \I__4755\ : Odrv4
    port map (
            O => \N__22436\,
            I => \uu2.w_addr_userZ0Z_4\
        );

    \I__4754\ : InMux
    port map (
            O => \N__22429\,
            I => \N__22416\
        );

    \I__4753\ : InMux
    port map (
            O => \N__22428\,
            I => \N__22416\
        );

    \I__4752\ : InMux
    port map (
            O => \N__22427\,
            I => \N__22416\
        );

    \I__4751\ : InMux
    port map (
            O => \N__22426\,
            I => \N__22409\
        );

    \I__4750\ : InMux
    port map (
            O => \N__22425\,
            I => \N__22409\
        );

    \I__4749\ : InMux
    port map (
            O => \N__22424\,
            I => \N__22409\
        );

    \I__4748\ : InMux
    port map (
            O => \N__22423\,
            I => \N__22406\
        );

    \I__4747\ : LocalMux
    port map (
            O => \N__22416\,
            I => \uu2.un28_w_addr_user_i\
        );

    \I__4746\ : LocalMux
    port map (
            O => \N__22409\,
            I => \uu2.un28_w_addr_user_i\
        );

    \I__4745\ : LocalMux
    port map (
            O => \N__22406\,
            I => \uu2.un28_w_addr_user_i\
        );

    \I__4744\ : InMux
    port map (
            O => \N__22399\,
            I => \N__22390\
        );

    \I__4743\ : InMux
    port map (
            O => \N__22398\,
            I => \N__22390\
        );

    \I__4742\ : InMux
    port map (
            O => \N__22397\,
            I => \N__22383\
        );

    \I__4741\ : InMux
    port map (
            O => \N__22396\,
            I => \N__22383\
        );

    \I__4740\ : InMux
    port map (
            O => \N__22395\,
            I => \N__22383\
        );

    \I__4739\ : LocalMux
    port map (
            O => \N__22390\,
            I => \uu2.un404_ci\
        );

    \I__4738\ : LocalMux
    port map (
            O => \N__22383\,
            I => \uu2.un404_ci\
        );

    \I__4737\ : CascadeMux
    port map (
            O => \N__22378\,
            I => \N__22375\
        );

    \I__4736\ : InMux
    port map (
            O => \N__22375\,
            I => \N__22371\
        );

    \I__4735\ : CascadeMux
    port map (
            O => \N__22374\,
            I => \N__22367\
        );

    \I__4734\ : LocalMux
    port map (
            O => \N__22371\,
            I => \N__22364\
        );

    \I__4733\ : InMux
    port map (
            O => \N__22370\,
            I => \N__22359\
        );

    \I__4732\ : InMux
    port map (
            O => \N__22367\,
            I => \N__22359\
        );

    \I__4731\ : Odrv4
    port map (
            O => \N__22364\,
            I => \uu2.un426_ci_3\
        );

    \I__4730\ : LocalMux
    port map (
            O => \N__22359\,
            I => \uu2.un426_ci_3\
        );

    \I__4729\ : InMux
    port map (
            O => \N__22354\,
            I => \N__22343\
        );

    \I__4728\ : InMux
    port map (
            O => \N__22353\,
            I => \N__22343\
        );

    \I__4727\ : InMux
    port map (
            O => \N__22352\,
            I => \N__22343\
        );

    \I__4726\ : InMux
    port map (
            O => \N__22351\,
            I => \N__22340\
        );

    \I__4725\ : InMux
    port map (
            O => \N__22350\,
            I => \N__22337\
        );

    \I__4724\ : LocalMux
    port map (
            O => \N__22343\,
            I => \N__22332\
        );

    \I__4723\ : LocalMux
    port map (
            O => \N__22340\,
            I => \N__22332\
        );

    \I__4722\ : LocalMux
    port map (
            O => \N__22337\,
            I => \uu2.w_addr_userZ0Z_6\
        );

    \I__4721\ : Odrv4
    port map (
            O => \N__22332\,
            I => \uu2.w_addr_userZ0Z_6\
        );

    \I__4720\ : SRMux
    port map (
            O => \N__22327\,
            I => \N__22323\
        );

    \I__4719\ : SRMux
    port map (
            O => \N__22326\,
            I => \N__22319\
        );

    \I__4718\ : LocalMux
    port map (
            O => \N__22323\,
            I => \N__22316\
        );

    \I__4717\ : SRMux
    port map (
            O => \N__22322\,
            I => \N__22313\
        );

    \I__4716\ : LocalMux
    port map (
            O => \N__22319\,
            I => \N__22307\
        );

    \I__4715\ : Span4Mux_h
    port map (
            O => \N__22316\,
            I => \N__22307\
        );

    \I__4714\ : LocalMux
    port map (
            O => \N__22313\,
            I => \N__22304\
        );

    \I__4713\ : InMux
    port map (
            O => \N__22312\,
            I => \N__22301\
        );

    \I__4712\ : Odrv4
    port map (
            O => \N__22307\,
            I => \uu2.w_addr_user_RNIMJ3O2Z0Z_2\
        );

    \I__4711\ : Odrv4
    port map (
            O => \N__22304\,
            I => \uu2.w_addr_user_RNIMJ3O2Z0Z_2\
        );

    \I__4710\ : LocalMux
    port map (
            O => \N__22301\,
            I => \uu2.w_addr_user_RNIMJ3O2Z0Z_2\
        );

    \I__4709\ : InMux
    port map (
            O => \N__22294\,
            I => \N__22285\
        );

    \I__4708\ : InMux
    port map (
            O => \N__22293\,
            I => \N__22285\
        );

    \I__4707\ : InMux
    port map (
            O => \N__22292\,
            I => \N__22285\
        );

    \I__4706\ : LocalMux
    port map (
            O => \N__22285\,
            I => \L3_tx_data_rdy\
        );

    \I__4705\ : CascadeMux
    port map (
            O => \N__22282\,
            I => \N__22277\
        );

    \I__4704\ : InMux
    port map (
            O => \N__22281\,
            I => \N__22272\
        );

    \I__4703\ : InMux
    port map (
            O => \N__22280\,
            I => \N__22272\
        );

    \I__4702\ : InMux
    port map (
            O => \N__22277\,
            I => \N__22269\
        );

    \I__4701\ : LocalMux
    port map (
            O => \N__22272\,
            I => \L3_tx_data_6\
        );

    \I__4700\ : LocalMux
    port map (
            O => \N__22269\,
            I => \L3_tx_data_6\
        );

    \I__4699\ : InMux
    port map (
            O => \N__22264\,
            I => \N__22261\
        );

    \I__4698\ : LocalMux
    port map (
            O => \N__22261\,
            I => \N__22256\
        );

    \I__4697\ : InMux
    port map (
            O => \N__22260\,
            I => \N__22251\
        );

    \I__4696\ : InMux
    port map (
            O => \N__22259\,
            I => \N__22251\
        );

    \I__4695\ : Span4Mux_h
    port map (
            O => \N__22256\,
            I => \N__22248\
        );

    \I__4694\ : LocalMux
    port map (
            O => \N__22251\,
            I => \Lab_UT.uu0.l_countZ0Z_3\
        );

    \I__4693\ : Odrv4
    port map (
            O => \N__22248\,
            I => \Lab_UT.uu0.l_countZ0Z_3\
        );

    \I__4692\ : InMux
    port map (
            O => \N__22243\,
            I => \N__22236\
        );

    \I__4691\ : InMux
    port map (
            O => \N__22242\,
            I => \N__22236\
        );

    \I__4690\ : InMux
    port map (
            O => \N__22241\,
            I => \N__22232\
        );

    \I__4689\ : LocalMux
    port map (
            O => \N__22236\,
            I => \N__22229\
        );

    \I__4688\ : InMux
    port map (
            O => \N__22235\,
            I => \N__22226\
        );

    \I__4687\ : LocalMux
    port map (
            O => \N__22232\,
            I => \Lab_UT.uu0.l_countZ0Z_2\
        );

    \I__4686\ : Odrv4
    port map (
            O => \N__22229\,
            I => \Lab_UT.uu0.l_countZ0Z_2\
        );

    \I__4685\ : LocalMux
    port map (
            O => \N__22226\,
            I => \Lab_UT.uu0.l_countZ0Z_2\
        );

    \I__4684\ : CascadeMux
    port map (
            O => \N__22219\,
            I => \Lab_UT.uu0.un66_ci_cascade_\
        );

    \I__4683\ : InMux
    port map (
            O => \N__22216\,
            I => \N__22208\
        );

    \I__4682\ : InMux
    port map (
            O => \N__22215\,
            I => \N__22208\
        );

    \I__4681\ : InMux
    port map (
            O => \N__22214\,
            I => \N__22205\
        );

    \I__4680\ : InMux
    port map (
            O => \N__22213\,
            I => \N__22202\
        );

    \I__4679\ : LocalMux
    port map (
            O => \N__22208\,
            I => \Lab_UT.uu0.l_countZ0Z_4\
        );

    \I__4678\ : LocalMux
    port map (
            O => \N__22205\,
            I => \Lab_UT.uu0.l_countZ0Z_4\
        );

    \I__4677\ : LocalMux
    port map (
            O => \N__22202\,
            I => \Lab_UT.uu0.l_countZ0Z_4\
        );

    \I__4676\ : InMux
    port map (
            O => \N__22195\,
            I => \N__22187\
        );

    \I__4675\ : InMux
    port map (
            O => \N__22194\,
            I => \N__22187\
        );

    \I__4674\ : InMux
    port map (
            O => \N__22193\,
            I => \N__22184\
        );

    \I__4673\ : InMux
    port map (
            O => \N__22192\,
            I => \N__22181\
        );

    \I__4672\ : LocalMux
    port map (
            O => \N__22187\,
            I => \Lab_UT.uu0.un66_ci\
        );

    \I__4671\ : LocalMux
    port map (
            O => \N__22184\,
            I => \Lab_UT.uu0.un66_ci\
        );

    \I__4670\ : LocalMux
    port map (
            O => \N__22181\,
            I => \Lab_UT.uu0.un66_ci\
        );

    \I__4669\ : CEMux
    port map (
            O => \N__22174\,
            I => \N__22159\
        );

    \I__4668\ : CEMux
    port map (
            O => \N__22173\,
            I => \N__22159\
        );

    \I__4667\ : CEMux
    port map (
            O => \N__22172\,
            I => \N__22159\
        );

    \I__4666\ : CEMux
    port map (
            O => \N__22171\,
            I => \N__22159\
        );

    \I__4665\ : CEMux
    port map (
            O => \N__22170\,
            I => \N__22159\
        );

    \I__4664\ : GlobalMux
    port map (
            O => \N__22159\,
            I => \N__22156\
        );

    \I__4663\ : gio2CtrlBuf
    port map (
            O => \N__22156\,
            I => \Lab_UT.uu0.un11_l_count_i_g\
        );

    \I__4662\ : InMux
    port map (
            O => \N__22153\,
            I => \N__22150\
        );

    \I__4661\ : LocalMux
    port map (
            O => \N__22150\,
            I => \N__22147\
        );

    \I__4660\ : Span4Mux_v
    port map (
            O => \N__22147\,
            I => \N__22143\
        );

    \I__4659\ : InMux
    port map (
            O => \N__22146\,
            I => \N__22140\
        );

    \I__4658\ : Span4Mux_h
    port map (
            O => \N__22143\,
            I => \N__22135\
        );

    \I__4657\ : LocalMux
    port map (
            O => \N__22140\,
            I => \N__22135\
        );

    \I__4656\ : Span4Mux_v
    port map (
            O => \N__22135\,
            I => \N__22132\
        );

    \I__4655\ : Odrv4
    port map (
            O => \N__22132\,
            I => \Lab_UT.uu0.delay_lineZ0Z_0\
        );

    \I__4654\ : InMux
    port map (
            O => \N__22129\,
            I => \N__22124\
        );

    \I__4653\ : InMux
    port map (
            O => \N__22128\,
            I => \N__22121\
        );

    \I__4652\ : InMux
    port map (
            O => \N__22127\,
            I => \N__22118\
        );

    \I__4651\ : LocalMux
    port map (
            O => \N__22124\,
            I => \Lab_UT.uu0.l_countZ0Z_5\
        );

    \I__4650\ : LocalMux
    port map (
            O => \N__22121\,
            I => \Lab_UT.uu0.l_countZ0Z_5\
        );

    \I__4649\ : LocalMux
    port map (
            O => \N__22118\,
            I => \Lab_UT.uu0.l_countZ0Z_5\
        );

    \I__4648\ : CascadeMux
    port map (
            O => \N__22111\,
            I => \N__22106\
        );

    \I__4647\ : CascadeMux
    port map (
            O => \N__22110\,
            I => \N__22103\
        );

    \I__4646\ : InMux
    port map (
            O => \N__22109\,
            I => \N__22096\
        );

    \I__4645\ : InMux
    port map (
            O => \N__22106\,
            I => \N__22096\
        );

    \I__4644\ : InMux
    port map (
            O => \N__22103\,
            I => \N__22096\
        );

    \I__4643\ : LocalMux
    port map (
            O => \N__22096\,
            I => \Lab_UT.uu0.l_precountZ0Z_3\
        );

    \I__4642\ : InMux
    port map (
            O => \N__22093\,
            I => \N__22083\
        );

    \I__4641\ : InMux
    port map (
            O => \N__22092\,
            I => \N__22083\
        );

    \I__4640\ : InMux
    port map (
            O => \N__22091\,
            I => \N__22083\
        );

    \I__4639\ : InMux
    port map (
            O => \N__22090\,
            I => \N__22080\
        );

    \I__4638\ : LocalMux
    port map (
            O => \N__22083\,
            I => \Lab_UT.uu0.l_countZ0Z_1\
        );

    \I__4637\ : LocalMux
    port map (
            O => \N__22080\,
            I => \Lab_UT.uu0.l_countZ0Z_1\
        );

    \I__4636\ : InMux
    port map (
            O => \N__22075\,
            I => \N__22072\
        );

    \I__4635\ : LocalMux
    port map (
            O => \N__22072\,
            I => \N__22068\
        );

    \I__4634\ : InMux
    port map (
            O => \N__22071\,
            I => \N__22065\
        );

    \I__4633\ : Span4Mux_h
    port map (
            O => \N__22068\,
            I => \N__22062\
        );

    \I__4632\ : LocalMux
    port map (
            O => \N__22065\,
            I => \Lab_UT.uu0.l_countZ0Z_18\
        );

    \I__4631\ : Odrv4
    port map (
            O => \N__22062\,
            I => \Lab_UT.uu0.l_countZ0Z_18\
        );

    \I__4630\ : InMux
    port map (
            O => \N__22057\,
            I => \N__22052\
        );

    \I__4629\ : InMux
    port map (
            O => \N__22056\,
            I => \N__22049\
        );

    \I__4628\ : InMux
    port map (
            O => \N__22055\,
            I => \N__22046\
        );

    \I__4627\ : LocalMux
    port map (
            O => \N__22052\,
            I => \Lab_UT.uu0.l_countZ0Z_15\
        );

    \I__4626\ : LocalMux
    port map (
            O => \N__22049\,
            I => \Lab_UT.uu0.l_countZ0Z_15\
        );

    \I__4625\ : LocalMux
    port map (
            O => \N__22046\,
            I => \Lab_UT.uu0.l_countZ0Z_15\
        );

    \I__4624\ : CascadeMux
    port map (
            O => \N__22039\,
            I => \Lab_UT.uu0.un4_l_count_11_cascade_\
        );

    \I__4623\ : InMux
    port map (
            O => \N__22036\,
            I => \N__22026\
        );

    \I__4622\ : InMux
    port map (
            O => \N__22035\,
            I => \N__22026\
        );

    \I__4621\ : InMux
    port map (
            O => \N__22034\,
            I => \N__22026\
        );

    \I__4620\ : InMux
    port map (
            O => \N__22033\,
            I => \N__22023\
        );

    \I__4619\ : LocalMux
    port map (
            O => \N__22026\,
            I => \Lab_UT.uu0.l_countZ0Z_6\
        );

    \I__4618\ : LocalMux
    port map (
            O => \N__22023\,
            I => \Lab_UT.uu0.l_countZ0Z_6\
        );

    \I__4617\ : InMux
    port map (
            O => \N__22018\,
            I => \N__22015\
        );

    \I__4616\ : LocalMux
    port map (
            O => \N__22015\,
            I => \N__22012\
        );

    \I__4615\ : Odrv4
    port map (
            O => \N__22012\,
            I => \Lab_UT.uu0.un4_l_count_12\
        );

    \I__4614\ : CascadeMux
    port map (
            O => \N__22009\,
            I => \Lab_UT.uu0.un4_l_count_16_cascade_\
        );

    \I__4613\ : InMux
    port map (
            O => \N__22006\,
            I => \N__22003\
        );

    \I__4612\ : LocalMux
    port map (
            O => \N__22003\,
            I => \Lab_UT.uu0.un4_l_count_18\
        );

    \I__4611\ : InMux
    port map (
            O => \N__22000\,
            I => \N__21996\
        );

    \I__4610\ : CascadeMux
    port map (
            O => \N__21999\,
            I => \N__21992\
        );

    \I__4609\ : LocalMux
    port map (
            O => \N__21996\,
            I => \N__21988\
        );

    \I__4608\ : CascadeMux
    port map (
            O => \N__21995\,
            I => \N__21983\
        );

    \I__4607\ : InMux
    port map (
            O => \N__21992\,
            I => \N__21980\
        );

    \I__4606\ : CascadeMux
    port map (
            O => \N__21991\,
            I => \N__21977\
        );

    \I__4605\ : Span4Mux_v
    port map (
            O => \N__21988\,
            I => \N__21974\
        );

    \I__4604\ : CascadeMux
    port map (
            O => \N__21987\,
            I => \N__21971\
        );

    \I__4603\ : InMux
    port map (
            O => \N__21986\,
            I => \N__21966\
        );

    \I__4602\ : InMux
    port map (
            O => \N__21983\,
            I => \N__21966\
        );

    \I__4601\ : LocalMux
    port map (
            O => \N__21980\,
            I => \N__21963\
        );

    \I__4600\ : InMux
    port map (
            O => \N__21977\,
            I => \N__21960\
        );

    \I__4599\ : Span4Mux_h
    port map (
            O => \N__21974\,
            I => \N__21957\
        );

    \I__4598\ : InMux
    port map (
            O => \N__21971\,
            I => \N__21954\
        );

    \I__4597\ : LocalMux
    port map (
            O => \N__21966\,
            I => \N__21949\
        );

    \I__4596\ : Span4Mux_v
    port map (
            O => \N__21963\,
            I => \N__21949\
        );

    \I__4595\ : LocalMux
    port map (
            O => \N__21960\,
            I => \N__21946\
        );

    \I__4594\ : Odrv4
    port map (
            O => \N__21957\,
            I => bu_rx_data_6_rep1
        );

    \I__4593\ : LocalMux
    port map (
            O => \N__21954\,
            I => bu_rx_data_6_rep1
        );

    \I__4592\ : Odrv4
    port map (
            O => \N__21949\,
            I => bu_rx_data_6_rep1
        );

    \I__4591\ : Odrv4
    port map (
            O => \N__21946\,
            I => bu_rx_data_6_rep1
        );

    \I__4590\ : InMux
    port map (
            O => \N__21937\,
            I => \N__21932\
        );

    \I__4589\ : InMux
    port map (
            O => \N__21936\,
            I => \N__21929\
        );

    \I__4588\ : InMux
    port map (
            O => \N__21935\,
            I => \N__21926\
        );

    \I__4587\ : LocalMux
    port map (
            O => \N__21932\,
            I => \N__21919\
        );

    \I__4586\ : LocalMux
    port map (
            O => \N__21929\,
            I => \N__21919\
        );

    \I__4585\ : LocalMux
    port map (
            O => \N__21926\,
            I => \N__21915\
        );

    \I__4584\ : InMux
    port map (
            O => \N__21925\,
            I => \N__21910\
        );

    \I__4583\ : InMux
    port map (
            O => \N__21924\,
            I => \N__21910\
        );

    \I__4582\ : Span4Mux_h
    port map (
            O => \N__21919\,
            I => \N__21907\
        );

    \I__4581\ : InMux
    port map (
            O => \N__21918\,
            I => \N__21904\
        );

    \I__4580\ : Odrv4
    port map (
            O => \N__21915\,
            I => bu_rx_data_5_rep1
        );

    \I__4579\ : LocalMux
    port map (
            O => \N__21910\,
            I => bu_rx_data_5_rep1
        );

    \I__4578\ : Odrv4
    port map (
            O => \N__21907\,
            I => bu_rx_data_5_rep1
        );

    \I__4577\ : LocalMux
    port map (
            O => \N__21904\,
            I => bu_rx_data_5_rep1
        );

    \I__4576\ : InMux
    port map (
            O => \N__21895\,
            I => \N__21892\
        );

    \I__4575\ : LocalMux
    port map (
            O => \N__21892\,
            I => \N__21888\
        );

    \I__4574\ : InMux
    port map (
            O => \N__21891\,
            I => \N__21885\
        );

    \I__4573\ : Span4Mux_h
    port map (
            O => \N__21888\,
            I => \N__21882\
        );

    \I__4572\ : LocalMux
    port map (
            O => \N__21885\,
            I => bu_rx_data_fast_3
        );

    \I__4571\ : Odrv4
    port map (
            O => \N__21882\,
            I => bu_rx_data_fast_3
        );

    \I__4570\ : InMux
    port map (
            O => \N__21877\,
            I => \N__21873\
        );

    \I__4569\ : InMux
    port map (
            O => \N__21876\,
            I => \N__21868\
        );

    \I__4568\ : LocalMux
    port map (
            O => \N__21873\,
            I => \N__21865\
        );

    \I__4567\ : InMux
    port map (
            O => \N__21872\,
            I => \N__21862\
        );

    \I__4566\ : InMux
    port map (
            O => \N__21871\,
            I => \N__21859\
        );

    \I__4565\ : LocalMux
    port map (
            O => \N__21868\,
            I => \N__21852\
        );

    \I__4564\ : Span4Mux_v
    port map (
            O => \N__21865\,
            I => \N__21852\
        );

    \I__4563\ : LocalMux
    port map (
            O => \N__21862\,
            I => \N__21852\
        );

    \I__4562\ : LocalMux
    port map (
            O => \N__21859\,
            I => \N__21849\
        );

    \I__4561\ : Span4Mux_h
    port map (
            O => \N__21852\,
            I => \N__21846\
        );

    \I__4560\ : Odrv12
    port map (
            O => \N__21849\,
            I => \buart.Z_rx.hhZ0Z_1\
        );

    \I__4559\ : Odrv4
    port map (
            O => \N__21846\,
            I => \buart.Z_rx.hhZ0Z_1\
        );

    \I__4558\ : InMux
    port map (
            O => \N__21841\,
            I => \N__21838\
        );

    \I__4557\ : LocalMux
    port map (
            O => \N__21838\,
            I => \N__21834\
        );

    \I__4556\ : InMux
    port map (
            O => \N__21837\,
            I => \N__21828\
        );

    \I__4555\ : Span4Mux_s3_h
    port map (
            O => \N__21834\,
            I => \N__21825\
        );

    \I__4554\ : InMux
    port map (
            O => \N__21833\,
            I => \N__21820\
        );

    \I__4553\ : InMux
    port map (
            O => \N__21832\,
            I => \N__21820\
        );

    \I__4552\ : CascadeMux
    port map (
            O => \N__21831\,
            I => \N__21816\
        );

    \I__4551\ : LocalMux
    port map (
            O => \N__21828\,
            I => \N__21813\
        );

    \I__4550\ : Span4Mux_h
    port map (
            O => \N__21825\,
            I => \N__21810\
        );

    \I__4549\ : LocalMux
    port map (
            O => \N__21820\,
            I => \N__21807\
        );

    \I__4548\ : InMux
    port map (
            O => \N__21819\,
            I => \N__21802\
        );

    \I__4547\ : InMux
    port map (
            O => \N__21816\,
            I => \N__21802\
        );

    \I__4546\ : Odrv4
    port map (
            O => \N__21813\,
            I => bu_rx_data_7_rep1
        );

    \I__4545\ : Odrv4
    port map (
            O => \N__21810\,
            I => bu_rx_data_7_rep1
        );

    \I__4544\ : Odrv4
    port map (
            O => \N__21807\,
            I => bu_rx_data_7_rep1
        );

    \I__4543\ : LocalMux
    port map (
            O => \N__21802\,
            I => bu_rx_data_7_rep1
        );

    \I__4542\ : InMux
    port map (
            O => \N__21793\,
            I => \N__21790\
        );

    \I__4541\ : LocalMux
    port map (
            O => \N__21790\,
            I => \N__21787\
        );

    \I__4540\ : Odrv4
    port map (
            O => \N__21787\,
            I => \Lab_UT.uu0.un44_ci\
        );

    \I__4539\ : CascadeMux
    port map (
            O => \N__21784\,
            I => \Lab_UT.uu0.un44_ci_cascade_\
        );

    \I__4538\ : CascadeMux
    port map (
            O => \N__21781\,
            I => \N__21777\
        );

    \I__4537\ : CascadeMux
    port map (
            O => \N__21780\,
            I => \N__21774\
        );

    \I__4536\ : InMux
    port map (
            O => \N__21777\,
            I => \N__21771\
        );

    \I__4535\ : InMux
    port map (
            O => \N__21774\,
            I => \N__21768\
        );

    \I__4534\ : LocalMux
    port map (
            O => \N__21771\,
            I => \N__21760\
        );

    \I__4533\ : LocalMux
    port map (
            O => \N__21768\,
            I => \N__21757\
        );

    \I__4532\ : CascadeMux
    port map (
            O => \N__21767\,
            I => \N__21753\
        );

    \I__4531\ : CascadeMux
    port map (
            O => \N__21766\,
            I => \N__21750\
        );

    \I__4530\ : InMux
    port map (
            O => \N__21765\,
            I => \N__21742\
        );

    \I__4529\ : InMux
    port map (
            O => \N__21764\,
            I => \N__21742\
        );

    \I__4528\ : InMux
    port map (
            O => \N__21763\,
            I => \N__21742\
        );

    \I__4527\ : Span4Mux_h
    port map (
            O => \N__21760\,
            I => \N__21739\
        );

    \I__4526\ : Span4Mux_h
    port map (
            O => \N__21757\,
            I => \N__21736\
        );

    \I__4525\ : InMux
    port map (
            O => \N__21756\,
            I => \N__21727\
        );

    \I__4524\ : InMux
    port map (
            O => \N__21753\,
            I => \N__21727\
        );

    \I__4523\ : InMux
    port map (
            O => \N__21750\,
            I => \N__21727\
        );

    \I__4522\ : InMux
    port map (
            O => \N__21749\,
            I => \N__21727\
        );

    \I__4521\ : LocalMux
    port map (
            O => \N__21742\,
            I => bu_rx_data_3_rep1
        );

    \I__4520\ : Odrv4
    port map (
            O => \N__21739\,
            I => bu_rx_data_3_rep1
        );

    \I__4519\ : Odrv4
    port map (
            O => \N__21736\,
            I => bu_rx_data_3_rep1
        );

    \I__4518\ : LocalMux
    port map (
            O => \N__21727\,
            I => bu_rx_data_3_rep1
        );

    \I__4517\ : CascadeMux
    port map (
            O => \N__21718\,
            I => \Lab_UT.dictrl.g1_5_1_cascade_\
        );

    \I__4516\ : InMux
    port map (
            O => \N__21715\,
            I => \N__21712\
        );

    \I__4515\ : LocalMux
    port map (
            O => \N__21712\,
            I => \N__21709\
        );

    \I__4514\ : Span4Mux_v
    port map (
            O => \N__21709\,
            I => \N__21706\
        );

    \I__4513\ : Odrv4
    port map (
            O => \N__21706\,
            I => \Lab_UT.dictrl.g1_7_1\
        );

    \I__4512\ : InMux
    port map (
            O => \N__21703\,
            I => \N__21700\
        );

    \I__4511\ : LocalMux
    port map (
            O => \N__21700\,
            I => \N__21692\
        );

    \I__4510\ : InMux
    port map (
            O => \N__21699\,
            I => \N__21689\
        );

    \I__4509\ : CascadeMux
    port map (
            O => \N__21698\,
            I => \N__21686\
        );

    \I__4508\ : InMux
    port map (
            O => \N__21697\,
            I => \N__21680\
        );

    \I__4507\ : InMux
    port map (
            O => \N__21696\,
            I => \N__21675\
        );

    \I__4506\ : InMux
    port map (
            O => \N__21695\,
            I => \N__21675\
        );

    \I__4505\ : Span4Mux_h
    port map (
            O => \N__21692\,
            I => \N__21672\
        );

    \I__4504\ : LocalMux
    port map (
            O => \N__21689\,
            I => \N__21669\
        );

    \I__4503\ : InMux
    port map (
            O => \N__21686\,
            I => \N__21660\
        );

    \I__4502\ : InMux
    port map (
            O => \N__21685\,
            I => \N__21660\
        );

    \I__4501\ : InMux
    port map (
            O => \N__21684\,
            I => \N__21660\
        );

    \I__4500\ : InMux
    port map (
            O => \N__21683\,
            I => \N__21660\
        );

    \I__4499\ : LocalMux
    port map (
            O => \N__21680\,
            I => bu_rx_data_2_rep1
        );

    \I__4498\ : LocalMux
    port map (
            O => \N__21675\,
            I => bu_rx_data_2_rep1
        );

    \I__4497\ : Odrv4
    port map (
            O => \N__21672\,
            I => bu_rx_data_2_rep1
        );

    \I__4496\ : Odrv12
    port map (
            O => \N__21669\,
            I => bu_rx_data_2_rep1
        );

    \I__4495\ : LocalMux
    port map (
            O => \N__21660\,
            I => bu_rx_data_2_rep1
        );

    \I__4494\ : InMux
    port map (
            O => \N__21649\,
            I => \N__21646\
        );

    \I__4493\ : LocalMux
    port map (
            O => \N__21646\,
            I => \N__21643\
        );

    \I__4492\ : Odrv4
    port map (
            O => \N__21643\,
            I => \Lab_UT.dictrl.g1_4_1\
        );

    \I__4491\ : InMux
    port map (
            O => \N__21640\,
            I => \N__21637\
        );

    \I__4490\ : LocalMux
    port map (
            O => \N__21637\,
            I => \Lab_UT.dictrl.currState_fast_3\
        );

    \I__4489\ : InMux
    port map (
            O => \N__21634\,
            I => \N__21631\
        );

    \I__4488\ : LocalMux
    port map (
            O => \N__21631\,
            I => \N__21628\
        );

    \I__4487\ : Odrv4
    port map (
            O => \N__21628\,
            I => \buart.Z_rx.G_30_0_o3_1_4\
        );

    \I__4486\ : InMux
    port map (
            O => \N__21625\,
            I => \N__21611\
        );

    \I__4485\ : InMux
    port map (
            O => \N__21624\,
            I => \N__21603\
        );

    \I__4484\ : InMux
    port map (
            O => \N__21623\,
            I => \N__21598\
        );

    \I__4483\ : InMux
    port map (
            O => \N__21622\,
            I => \N__21598\
        );

    \I__4482\ : InMux
    port map (
            O => \N__21621\,
            I => \N__21581\
        );

    \I__4481\ : InMux
    port map (
            O => \N__21620\,
            I => \N__21581\
        );

    \I__4480\ : InMux
    port map (
            O => \N__21619\,
            I => \N__21581\
        );

    \I__4479\ : InMux
    port map (
            O => \N__21618\,
            I => \N__21581\
        );

    \I__4478\ : InMux
    port map (
            O => \N__21617\,
            I => \N__21581\
        );

    \I__4477\ : InMux
    port map (
            O => \N__21616\,
            I => \N__21581\
        );

    \I__4476\ : InMux
    port map (
            O => \N__21615\,
            I => \N__21581\
        );

    \I__4475\ : InMux
    port map (
            O => \N__21614\,
            I => \N__21581\
        );

    \I__4474\ : LocalMux
    port map (
            O => \N__21611\,
            I => \N__21578\
        );

    \I__4473\ : CascadeMux
    port map (
            O => \N__21610\,
            I => \N__21569\
        );

    \I__4472\ : CascadeMux
    port map (
            O => \N__21609\,
            I => \N__21565\
        );

    \I__4471\ : InMux
    port map (
            O => \N__21608\,
            I => \N__21562\
        );

    \I__4470\ : InMux
    port map (
            O => \N__21607\,
            I => \N__21559\
        );

    \I__4469\ : InMux
    port map (
            O => \N__21606\,
            I => \N__21556\
        );

    \I__4468\ : LocalMux
    port map (
            O => \N__21603\,
            I => \N__21553\
        );

    \I__4467\ : LocalMux
    port map (
            O => \N__21598\,
            I => \N__21550\
        );

    \I__4466\ : LocalMux
    port map (
            O => \N__21581\,
            I => \N__21547\
        );

    \I__4465\ : Span4Mux_s1_h
    port map (
            O => \N__21578\,
            I => \N__21544\
        );

    \I__4464\ : InMux
    port map (
            O => \N__21577\,
            I => \N__21537\
        );

    \I__4463\ : InMux
    port map (
            O => \N__21576\,
            I => \N__21537\
        );

    \I__4462\ : InMux
    port map (
            O => \N__21575\,
            I => \N__21537\
        );

    \I__4461\ : InMux
    port map (
            O => \N__21574\,
            I => \N__21529\
        );

    \I__4460\ : InMux
    port map (
            O => \N__21573\,
            I => \N__21529\
        );

    \I__4459\ : InMux
    port map (
            O => \N__21572\,
            I => \N__21529\
        );

    \I__4458\ : InMux
    port map (
            O => \N__21569\,
            I => \N__21522\
        );

    \I__4457\ : InMux
    port map (
            O => \N__21568\,
            I => \N__21522\
        );

    \I__4456\ : InMux
    port map (
            O => \N__21565\,
            I => \N__21522\
        );

    \I__4455\ : LocalMux
    port map (
            O => \N__21562\,
            I => \N__21508\
        );

    \I__4454\ : LocalMux
    port map (
            O => \N__21559\,
            I => \N__21508\
        );

    \I__4453\ : LocalMux
    port map (
            O => \N__21556\,
            I => \N__21501\
        );

    \I__4452\ : Span4Mux_v
    port map (
            O => \N__21553\,
            I => \N__21501\
        );

    \I__4451\ : Span4Mux_v
    port map (
            O => \N__21550\,
            I => \N__21501\
        );

    \I__4450\ : Span4Mux_h
    port map (
            O => \N__21547\,
            I => \N__21496\
        );

    \I__4449\ : Span4Mux_h
    port map (
            O => \N__21544\,
            I => \N__21496\
        );

    \I__4448\ : LocalMux
    port map (
            O => \N__21537\,
            I => \N__21493\
        );

    \I__4447\ : InMux
    port map (
            O => \N__21536\,
            I => \N__21490\
        );

    \I__4446\ : LocalMux
    port map (
            O => \N__21529\,
            I => \N__21485\
        );

    \I__4445\ : LocalMux
    port map (
            O => \N__21522\,
            I => \N__21485\
        );

    \I__4444\ : InMux
    port map (
            O => \N__21521\,
            I => \N__21470\
        );

    \I__4443\ : InMux
    port map (
            O => \N__21520\,
            I => \N__21470\
        );

    \I__4442\ : InMux
    port map (
            O => \N__21519\,
            I => \N__21470\
        );

    \I__4441\ : InMux
    port map (
            O => \N__21518\,
            I => \N__21470\
        );

    \I__4440\ : InMux
    port map (
            O => \N__21517\,
            I => \N__21470\
        );

    \I__4439\ : InMux
    port map (
            O => \N__21516\,
            I => \N__21470\
        );

    \I__4438\ : InMux
    port map (
            O => \N__21515\,
            I => \N__21470\
        );

    \I__4437\ : InMux
    port map (
            O => \N__21514\,
            I => \N__21465\
        );

    \I__4436\ : InMux
    port map (
            O => \N__21513\,
            I => \N__21465\
        );

    \I__4435\ : Span4Mux_v
    port map (
            O => \N__21508\,
            I => \N__21462\
        );

    \I__4434\ : Odrv4
    port map (
            O => \N__21501\,
            I => \Lab_UT.dictrl.nextStateZ0Z_3\
        );

    \I__4433\ : Odrv4
    port map (
            O => \N__21496\,
            I => \Lab_UT.dictrl.nextStateZ0Z_3\
        );

    \I__4432\ : Odrv12
    port map (
            O => \N__21493\,
            I => \Lab_UT.dictrl.nextStateZ0Z_3\
        );

    \I__4431\ : LocalMux
    port map (
            O => \N__21490\,
            I => \Lab_UT.dictrl.nextStateZ0Z_3\
        );

    \I__4430\ : Odrv4
    port map (
            O => \N__21485\,
            I => \Lab_UT.dictrl.nextStateZ0Z_3\
        );

    \I__4429\ : LocalMux
    port map (
            O => \N__21470\,
            I => \Lab_UT.dictrl.nextStateZ0Z_3\
        );

    \I__4428\ : LocalMux
    port map (
            O => \N__21465\,
            I => \Lab_UT.dictrl.nextStateZ0Z_3\
        );

    \I__4427\ : Odrv4
    port map (
            O => \N__21462\,
            I => \Lab_UT.dictrl.nextStateZ0Z_3\
        );

    \I__4426\ : InMux
    port map (
            O => \N__21445\,
            I => \N__21438\
        );

    \I__4425\ : InMux
    port map (
            O => \N__21444\,
            I => \N__21435\
        );

    \I__4424\ : InMux
    port map (
            O => \N__21443\,
            I => \N__21430\
        );

    \I__4423\ : InMux
    port map (
            O => \N__21442\,
            I => \N__21430\
        );

    \I__4422\ : InMux
    port map (
            O => \N__21441\,
            I => \N__21427\
        );

    \I__4421\ : LocalMux
    port map (
            O => \N__21438\,
            I => \N__21420\
        );

    \I__4420\ : LocalMux
    port map (
            O => \N__21435\,
            I => \N__21420\
        );

    \I__4419\ : LocalMux
    port map (
            O => \N__21430\,
            I => \N__21420\
        );

    \I__4418\ : LocalMux
    port map (
            O => \N__21427\,
            I => bu_rx_data_4_rep1
        );

    \I__4417\ : Odrv12
    port map (
            O => \N__21420\,
            I => bu_rx_data_4_rep1
        );

    \I__4416\ : InMux
    port map (
            O => \N__21415\,
            I => \N__21411\
        );

    \I__4415\ : InMux
    port map (
            O => \N__21414\,
            I => \N__21408\
        );

    \I__4414\ : LocalMux
    port map (
            O => \N__21411\,
            I => \N__21403\
        );

    \I__4413\ : LocalMux
    port map (
            O => \N__21408\,
            I => \N__21400\
        );

    \I__4412\ : InMux
    port map (
            O => \N__21407\,
            I => \N__21395\
        );

    \I__4411\ : InMux
    port map (
            O => \N__21406\,
            I => \N__21395\
        );

    \I__4410\ : Span4Mux_v
    port map (
            O => \N__21403\,
            I => \N__21384\
        );

    \I__4409\ : Span4Mux_s2_v
    port map (
            O => \N__21400\,
            I => \N__21384\
        );

    \I__4408\ : LocalMux
    port map (
            O => \N__21395\,
            I => \N__21381\
        );

    \I__4407\ : InMux
    port map (
            O => \N__21394\,
            I => \N__21376\
        );

    \I__4406\ : InMux
    port map (
            O => \N__21393\,
            I => \N__21376\
        );

    \I__4405\ : InMux
    port map (
            O => \N__21392\,
            I => \N__21367\
        );

    \I__4404\ : InMux
    port map (
            O => \N__21391\,
            I => \N__21367\
        );

    \I__4403\ : InMux
    port map (
            O => \N__21390\,
            I => \N__21367\
        );

    \I__4402\ : InMux
    port map (
            O => \N__21389\,
            I => \N__21367\
        );

    \I__4401\ : Odrv4
    port map (
            O => \N__21384\,
            I => bu_rx_data_1_rep1
        );

    \I__4400\ : Odrv12
    port map (
            O => \N__21381\,
            I => bu_rx_data_1_rep1
        );

    \I__4399\ : LocalMux
    port map (
            O => \N__21376\,
            I => bu_rx_data_1_rep1
        );

    \I__4398\ : LocalMux
    port map (
            O => \N__21367\,
            I => bu_rx_data_1_rep1
        );

    \I__4397\ : InMux
    port map (
            O => \N__21358\,
            I => \N__21355\
        );

    \I__4396\ : LocalMux
    port map (
            O => \N__21355\,
            I => \Lab_UT.dictrl.decoder.g0Z0Z_3\
        );

    \I__4395\ : InMux
    port map (
            O => \N__21352\,
            I => \N__21348\
        );

    \I__4394\ : InMux
    port map (
            O => \N__21351\,
            I => \N__21343\
        );

    \I__4393\ : LocalMux
    port map (
            O => \N__21348\,
            I => \N__21340\
        );

    \I__4392\ : InMux
    port map (
            O => \N__21347\,
            I => \N__21335\
        );

    \I__4391\ : InMux
    port map (
            O => \N__21346\,
            I => \N__21335\
        );

    \I__4390\ : LocalMux
    port map (
            O => \N__21343\,
            I => \N__21330\
        );

    \I__4389\ : Span4Mux_v
    port map (
            O => \N__21340\,
            I => \N__21330\
        );

    \I__4388\ : LocalMux
    port map (
            O => \N__21335\,
            I => bu_rx_data_0_rep1
        );

    \I__4387\ : Odrv4
    port map (
            O => \N__21330\,
            I => bu_rx_data_0_rep1
        );

    \I__4386\ : InMux
    port map (
            O => \N__21325\,
            I => \N__21322\
        );

    \I__4385\ : LocalMux
    port map (
            O => \N__21322\,
            I => \Lab_UT.dictrl.r_dicLdMtens14_i_6\
        );

    \I__4384\ : InMux
    port map (
            O => \N__21319\,
            I => \N__21316\
        );

    \I__4383\ : LocalMux
    port map (
            O => \N__21316\,
            I => \N__21313\
        );

    \I__4382\ : Span4Mux_h
    port map (
            O => \N__21313\,
            I => \N__21310\
        );

    \I__4381\ : Odrv4
    port map (
            O => \N__21310\,
            I => \Lab_UT.dictrl.r_dicLdMtens20_i_6\
        );

    \I__4380\ : InMux
    port map (
            O => \N__21307\,
            I => \N__21304\
        );

    \I__4379\ : LocalMux
    port map (
            O => \N__21304\,
            I => \N__21301\
        );

    \I__4378\ : Span4Mux_h
    port map (
            O => \N__21301\,
            I => \N__21298\
        );

    \I__4377\ : Odrv4
    port map (
            O => \N__21298\,
            I => \Lab_UT.dictrl.r_enable3_3_iv_1\
        );

    \I__4376\ : CascadeMux
    port map (
            O => \N__21295\,
            I => \buart.Z_rx.G_30_0_o3_1_0_cascade_\
        );

    \I__4375\ : InMux
    port map (
            O => \N__21292\,
            I => \N__21287\
        );

    \I__4374\ : InMux
    port map (
            O => \N__21291\,
            I => \N__21281\
        );

    \I__4373\ : InMux
    port map (
            O => \N__21290\,
            I => \N__21281\
        );

    \I__4372\ : LocalMux
    port map (
            O => \N__21287\,
            I => \N__21278\
        );

    \I__4371\ : InMux
    port map (
            O => \N__21286\,
            I => \N__21275\
        );

    \I__4370\ : LocalMux
    port map (
            O => \N__21281\,
            I => \Lab_UT_dictrl_decoder_de_cr_1\
        );

    \I__4369\ : Odrv4
    port map (
            O => \N__21278\,
            I => \Lab_UT_dictrl_decoder_de_cr_1\
        );

    \I__4368\ : LocalMux
    port map (
            O => \N__21275\,
            I => \Lab_UT_dictrl_decoder_de_cr_1\
        );

    \I__4367\ : CascadeMux
    port map (
            O => \N__21268\,
            I => \N__21261\
        );

    \I__4366\ : InMux
    port map (
            O => \N__21267\,
            I => \N__21254\
        );

    \I__4365\ : InMux
    port map (
            O => \N__21266\,
            I => \N__21254\
        );

    \I__4364\ : CascadeMux
    port map (
            O => \N__21265\,
            I => \N__21251\
        );

    \I__4363\ : CascadeMux
    port map (
            O => \N__21264\,
            I => \N__21247\
        );

    \I__4362\ : InMux
    port map (
            O => \N__21261\,
            I => \N__21241\
        );

    \I__4361\ : InMux
    port map (
            O => \N__21260\,
            I => \N__21238\
        );

    \I__4360\ : InMux
    port map (
            O => \N__21259\,
            I => \N__21235\
        );

    \I__4359\ : LocalMux
    port map (
            O => \N__21254\,
            I => \N__21231\
        );

    \I__4358\ : InMux
    port map (
            O => \N__21251\,
            I => \N__21228\
        );

    \I__4357\ : InMux
    port map (
            O => \N__21250\,
            I => \N__21223\
        );

    \I__4356\ : InMux
    port map (
            O => \N__21247\,
            I => \N__21223\
        );

    \I__4355\ : InMux
    port map (
            O => \N__21246\,
            I => \N__21219\
        );

    \I__4354\ : InMux
    port map (
            O => \N__21245\,
            I => \N__21215\
        );

    \I__4353\ : CascadeMux
    port map (
            O => \N__21244\,
            I => \N__21212\
        );

    \I__4352\ : LocalMux
    port map (
            O => \N__21241\,
            I => \N__21207\
        );

    \I__4351\ : LocalMux
    port map (
            O => \N__21238\,
            I => \N__21207\
        );

    \I__4350\ : LocalMux
    port map (
            O => \N__21235\,
            I => \N__21204\
        );

    \I__4349\ : InMux
    port map (
            O => \N__21234\,
            I => \N__21201\
        );

    \I__4348\ : Span4Mux_v
    port map (
            O => \N__21231\,
            I => \N__21194\
        );

    \I__4347\ : LocalMux
    port map (
            O => \N__21228\,
            I => \N__21194\
        );

    \I__4346\ : LocalMux
    port map (
            O => \N__21223\,
            I => \N__21194\
        );

    \I__4345\ : InMux
    port map (
            O => \N__21222\,
            I => \N__21191\
        );

    \I__4344\ : LocalMux
    port map (
            O => \N__21219\,
            I => \N__21188\
        );

    \I__4343\ : InMux
    port map (
            O => \N__21218\,
            I => \N__21185\
        );

    \I__4342\ : LocalMux
    port map (
            O => \N__21215\,
            I => \N__21182\
        );

    \I__4341\ : InMux
    port map (
            O => \N__21212\,
            I => \N__21179\
        );

    \I__4340\ : Span4Mux_v
    port map (
            O => \N__21207\,
            I => \N__21176\
        );

    \I__4339\ : Span4Mux_h
    port map (
            O => \N__21204\,
            I => \N__21171\
        );

    \I__4338\ : LocalMux
    port map (
            O => \N__21201\,
            I => \N__21171\
        );

    \I__4337\ : Span4Mux_v
    port map (
            O => \N__21194\,
            I => \N__21168\
        );

    \I__4336\ : LocalMux
    port map (
            O => \N__21191\,
            I => \N__21165\
        );

    \I__4335\ : Span4Mux_v
    port map (
            O => \N__21188\,
            I => \N__21160\
        );

    \I__4334\ : LocalMux
    port map (
            O => \N__21185\,
            I => \N__21160\
        );

    \I__4333\ : Span4Mux_s3_h
    port map (
            O => \N__21182\,
            I => \N__21157\
        );

    \I__4332\ : LocalMux
    port map (
            O => \N__21179\,
            I => \N__21152\
        );

    \I__4331\ : Span4Mux_h
    port map (
            O => \N__21176\,
            I => \N__21152\
        );

    \I__4330\ : Span4Mux_v
    port map (
            O => \N__21171\,
            I => \N__21147\
        );

    \I__4329\ : Span4Mux_h
    port map (
            O => \N__21168\,
            I => \N__21147\
        );

    \I__4328\ : Odrv12
    port map (
            O => \N__21165\,
            I => \Lab_UT.dictrl.currStateZ0Z_0\
        );

    \I__4327\ : Odrv4
    port map (
            O => \N__21160\,
            I => \Lab_UT.dictrl.currStateZ0Z_0\
        );

    \I__4326\ : Odrv4
    port map (
            O => \N__21157\,
            I => \Lab_UT.dictrl.currStateZ0Z_0\
        );

    \I__4325\ : Odrv4
    port map (
            O => \N__21152\,
            I => \Lab_UT.dictrl.currStateZ0Z_0\
        );

    \I__4324\ : Odrv4
    port map (
            O => \N__21147\,
            I => \Lab_UT.dictrl.currStateZ0Z_0\
        );

    \I__4323\ : CascadeMux
    port map (
            O => \N__21136\,
            I => \N_6_cascade_\
        );

    \I__4322\ : InMux
    port map (
            O => \N__21133\,
            I => \N__21130\
        );

    \I__4321\ : LocalMux
    port map (
            O => \N__21130\,
            I => \N__21127\
        );

    \I__4320\ : Span4Mux_s3_h
    port map (
            O => \N__21127\,
            I => \N__21124\
        );

    \I__4319\ : Span4Mux_h
    port map (
            O => \N__21124\,
            I => \N__21121\
        );

    \I__4318\ : Odrv4
    port map (
            O => \N__21121\,
            I => \Lab_UT.dictrl.N_21_0\
        );

    \I__4317\ : InMux
    port map (
            O => \N__21118\,
            I => \N__21115\
        );

    \I__4316\ : LocalMux
    port map (
            O => \N__21115\,
            I => \resetGen.escKey_4_0\
        );

    \I__4315\ : InMux
    port map (
            O => \N__21112\,
            I => \N__21104\
        );

    \I__4314\ : InMux
    port map (
            O => \N__21111\,
            I => \N__21099\
        );

    \I__4313\ : InMux
    port map (
            O => \N__21110\,
            I => \N__21099\
        );

    \I__4312\ : InMux
    port map (
            O => \N__21109\,
            I => \N__21087\
        );

    \I__4311\ : InMux
    port map (
            O => \N__21108\,
            I => \N__21084\
        );

    \I__4310\ : InMux
    port map (
            O => \N__21107\,
            I => \N__21081\
        );

    \I__4309\ : LocalMux
    port map (
            O => \N__21104\,
            I => \N__21076\
        );

    \I__4308\ : LocalMux
    port map (
            O => \N__21099\,
            I => \N__21076\
        );

    \I__4307\ : InMux
    port map (
            O => \N__21098\,
            I => \N__21073\
        );

    \I__4306\ : InMux
    port map (
            O => \N__21097\,
            I => \N__21054\
        );

    \I__4305\ : InMux
    port map (
            O => \N__21096\,
            I => \N__21054\
        );

    \I__4304\ : InMux
    port map (
            O => \N__21095\,
            I => \N__21054\
        );

    \I__4303\ : InMux
    port map (
            O => \N__21094\,
            I => \N__21054\
        );

    \I__4302\ : InMux
    port map (
            O => \N__21093\,
            I => \N__21054\
        );

    \I__4301\ : InMux
    port map (
            O => \N__21092\,
            I => \N__21054\
        );

    \I__4300\ : InMux
    port map (
            O => \N__21091\,
            I => \N__21054\
        );

    \I__4299\ : InMux
    port map (
            O => \N__21090\,
            I => \N__21054\
        );

    \I__4298\ : LocalMux
    port map (
            O => \N__21087\,
            I => \N__21051\
        );

    \I__4297\ : LocalMux
    port map (
            O => \N__21084\,
            I => \N__21048\
        );

    \I__4296\ : LocalMux
    port map (
            O => \N__21081\,
            I => \N__21045\
        );

    \I__4295\ : Span4Mux_v
    port map (
            O => \N__21076\,
            I => \N__21023\
        );

    \I__4294\ : LocalMux
    port map (
            O => \N__21073\,
            I => \N__21023\
        );

    \I__4293\ : InMux
    port map (
            O => \N__21072\,
            I => \N__21020\
        );

    \I__4292\ : InMux
    port map (
            O => \N__21071\,
            I => \N__21017\
        );

    \I__4291\ : LocalMux
    port map (
            O => \N__21054\,
            I => \N__21008\
        );

    \I__4290\ : Span4Mux_h
    port map (
            O => \N__21051\,
            I => \N__21008\
        );

    \I__4289\ : Span4Mux_v
    port map (
            O => \N__21048\,
            I => \N__21008\
        );

    \I__4288\ : Span4Mux_v
    port map (
            O => \N__21045\,
            I => \N__21008\
        );

    \I__4287\ : InMux
    port map (
            O => \N__21044\,
            I => \N__21001\
        );

    \I__4286\ : InMux
    port map (
            O => \N__21043\,
            I => \N__21001\
        );

    \I__4285\ : InMux
    port map (
            O => \N__21042\,
            I => \N__21001\
        );

    \I__4284\ : InMux
    port map (
            O => \N__21041\,
            I => \N__20990\
        );

    \I__4283\ : InMux
    port map (
            O => \N__21040\,
            I => \N__20990\
        );

    \I__4282\ : InMux
    port map (
            O => \N__21039\,
            I => \N__20990\
        );

    \I__4281\ : InMux
    port map (
            O => \N__21038\,
            I => \N__20990\
        );

    \I__4280\ : InMux
    port map (
            O => \N__21037\,
            I => \N__20990\
        );

    \I__4279\ : InMux
    port map (
            O => \N__21036\,
            I => \N__20985\
        );

    \I__4278\ : InMux
    port map (
            O => \N__21035\,
            I => \N__20985\
        );

    \I__4277\ : InMux
    port map (
            O => \N__21034\,
            I => \N__20970\
        );

    \I__4276\ : InMux
    port map (
            O => \N__21033\,
            I => \N__20970\
        );

    \I__4275\ : InMux
    port map (
            O => \N__21032\,
            I => \N__20970\
        );

    \I__4274\ : InMux
    port map (
            O => \N__21031\,
            I => \N__20970\
        );

    \I__4273\ : InMux
    port map (
            O => \N__21030\,
            I => \N__20970\
        );

    \I__4272\ : InMux
    port map (
            O => \N__21029\,
            I => \N__20970\
        );

    \I__4271\ : InMux
    port map (
            O => \N__21028\,
            I => \N__20970\
        );

    \I__4270\ : Span4Mux_h
    port map (
            O => \N__21023\,
            I => \N__20967\
        );

    \I__4269\ : LocalMux
    port map (
            O => \N__21020\,
            I => \Lab_UT.dictrl.nextStateZ0Z_0\
        );

    \I__4268\ : LocalMux
    port map (
            O => \N__21017\,
            I => \Lab_UT.dictrl.nextStateZ0Z_0\
        );

    \I__4267\ : Odrv4
    port map (
            O => \N__21008\,
            I => \Lab_UT.dictrl.nextStateZ0Z_0\
        );

    \I__4266\ : LocalMux
    port map (
            O => \N__21001\,
            I => \Lab_UT.dictrl.nextStateZ0Z_0\
        );

    \I__4265\ : LocalMux
    port map (
            O => \N__20990\,
            I => \Lab_UT.dictrl.nextStateZ0Z_0\
        );

    \I__4264\ : LocalMux
    port map (
            O => \N__20985\,
            I => \Lab_UT.dictrl.nextStateZ0Z_0\
        );

    \I__4263\ : LocalMux
    port map (
            O => \N__20970\,
            I => \Lab_UT.dictrl.nextStateZ0Z_0\
        );

    \I__4262\ : Odrv4
    port map (
            O => \N__20967\,
            I => \Lab_UT.dictrl.nextStateZ0Z_0\
        );

    \I__4261\ : CascadeMux
    port map (
            O => \N__20950\,
            I => \N__20946\
        );

    \I__4260\ : InMux
    port map (
            O => \N__20949\,
            I => \N__20941\
        );

    \I__4259\ : InMux
    port map (
            O => \N__20946\,
            I => \N__20941\
        );

    \I__4258\ : LocalMux
    port map (
            O => \N__20941\,
            I => \N__20932\
        );

    \I__4257\ : CascadeMux
    port map (
            O => \N__20940\,
            I => \N__20929\
        );

    \I__4256\ : CascadeMux
    port map (
            O => \N__20939\,
            I => \N__20926\
        );

    \I__4255\ : InMux
    port map (
            O => \N__20938\,
            I => \N__20923\
        );

    \I__4254\ : InMux
    port map (
            O => \N__20937\,
            I => \N__20916\
        );

    \I__4253\ : InMux
    port map (
            O => \N__20936\,
            I => \N__20916\
        );

    \I__4252\ : InMux
    port map (
            O => \N__20935\,
            I => \N__20916\
        );

    \I__4251\ : Span4Mux_h
    port map (
            O => \N__20932\,
            I => \N__20913\
        );

    \I__4250\ : InMux
    port map (
            O => \N__20929\,
            I => \N__20910\
        );

    \I__4249\ : InMux
    port map (
            O => \N__20926\,
            I => \N__20907\
        );

    \I__4248\ : LocalMux
    port map (
            O => \N__20923\,
            I => \N__20904\
        );

    \I__4247\ : LocalMux
    port map (
            O => \N__20916\,
            I => \N__20901\
        );

    \I__4246\ : Span4Mux_v
    port map (
            O => \N__20913\,
            I => \N__20895\
        );

    \I__4245\ : LocalMux
    port map (
            O => \N__20910\,
            I => \N__20895\
        );

    \I__4244\ : LocalMux
    port map (
            O => \N__20907\,
            I => \N__20892\
        );

    \I__4243\ : Span4Mux_v
    port map (
            O => \N__20904\,
            I => \N__20886\
        );

    \I__4242\ : Span4Mux_h
    port map (
            O => \N__20901\,
            I => \N__20886\
        );

    \I__4241\ : InMux
    port map (
            O => \N__20900\,
            I => \N__20883\
        );

    \I__4240\ : Span4Mux_h
    port map (
            O => \N__20895\,
            I => \N__20880\
        );

    \I__4239\ : Span4Mux_h
    port map (
            O => \N__20892\,
            I => \N__20877\
        );

    \I__4238\ : InMux
    port map (
            O => \N__20891\,
            I => \N__20874\
        );

    \I__4237\ : Span4Mux_h
    port map (
            O => \N__20886\,
            I => \N__20871\
        );

    \I__4236\ : LocalMux
    port map (
            O => \N__20883\,
            I => \Lab_UT.dictrl.currState_0_rep2\
        );

    \I__4235\ : Odrv4
    port map (
            O => \N__20880\,
            I => \Lab_UT.dictrl.currState_0_rep2\
        );

    \I__4234\ : Odrv4
    port map (
            O => \N__20877\,
            I => \Lab_UT.dictrl.currState_0_rep2\
        );

    \I__4233\ : LocalMux
    port map (
            O => \N__20874\,
            I => \Lab_UT.dictrl.currState_0_rep2\
        );

    \I__4232\ : Odrv4
    port map (
            O => \N__20871\,
            I => \Lab_UT.dictrl.currState_0_rep2\
        );

    \I__4231\ : CascadeMux
    port map (
            O => \N__20860\,
            I => \Lab_UT.dictrl.g0_7_cascade_\
        );

    \I__4230\ : CascadeMux
    port map (
            O => \N__20857\,
            I => \N__20854\
        );

    \I__4229\ : InMux
    port map (
            O => \N__20854\,
            I => \N__20851\
        );

    \I__4228\ : LocalMux
    port map (
            O => \N__20851\,
            I => \N__20848\
        );

    \I__4227\ : Span4Mux_h
    port map (
            O => \N__20848\,
            I => \N__20845\
        );

    \I__4226\ : Span4Mux_v
    port map (
            O => \N__20845\,
            I => \N__20842\
        );

    \I__4225\ : Odrv4
    port map (
            O => \N__20842\,
            I => \Lab_UT.dictrl.g0_10\
        );

    \I__4224\ : InMux
    port map (
            O => \N__20839\,
            I => \N__20835\
        );

    \I__4223\ : InMux
    port map (
            O => \N__20838\,
            I => \N__20832\
        );

    \I__4222\ : LocalMux
    port map (
            O => \N__20835\,
            I => \N__20829\
        );

    \I__4221\ : LocalMux
    port map (
            O => \N__20832\,
            I => bu_rx_data_fast_1
        );

    \I__4220\ : Odrv4
    port map (
            O => \N__20829\,
            I => bu_rx_data_fast_1
        );

    \I__4219\ : InMux
    port map (
            O => \N__20824\,
            I => \N__20821\
        );

    \I__4218\ : LocalMux
    port map (
            O => \N__20821\,
            I => \N__20818\
        );

    \I__4217\ : Odrv12
    port map (
            O => \N__20818\,
            I => \Lab_UT.dictrl.r_dicLdMtens16\
        );

    \I__4216\ : CascadeMux
    port map (
            O => \N__20815\,
            I => \N__20802\
        );

    \I__4215\ : InMux
    port map (
            O => \N__20814\,
            I => \N__20799\
        );

    \I__4214\ : InMux
    port map (
            O => \N__20813\,
            I => \N__20796\
        );

    \I__4213\ : CascadeMux
    port map (
            O => \N__20812\,
            I => \N__20789\
        );

    \I__4212\ : CascadeMux
    port map (
            O => \N__20811\,
            I => \N__20786\
        );

    \I__4211\ : CascadeMux
    port map (
            O => \N__20810\,
            I => \N__20783\
        );

    \I__4210\ : CascadeMux
    port map (
            O => \N__20809\,
            I => \N__20780\
        );

    \I__4209\ : CascadeMux
    port map (
            O => \N__20808\,
            I => \N__20777\
        );

    \I__4208\ : CascadeMux
    port map (
            O => \N__20807\,
            I => \N__20774\
        );

    \I__4207\ : CascadeMux
    port map (
            O => \N__20806\,
            I => \N__20771\
        );

    \I__4206\ : CascadeMux
    port map (
            O => \N__20805\,
            I => \N__20768\
        );

    \I__4205\ : InMux
    port map (
            O => \N__20802\,
            I => \N__20764\
        );

    \I__4204\ : LocalMux
    port map (
            O => \N__20799\,
            I => \N__20761\
        );

    \I__4203\ : LocalMux
    port map (
            O => \N__20796\,
            I => \N__20758\
        );

    \I__4202\ : CascadeMux
    port map (
            O => \N__20795\,
            I => \N__20752\
        );

    \I__4201\ : CascadeMux
    port map (
            O => \N__20794\,
            I => \N__20748\
        );

    \I__4200\ : CascadeMux
    port map (
            O => \N__20793\,
            I => \N__20743\
        );

    \I__4199\ : CascadeMux
    port map (
            O => \N__20792\,
            I => \N__20739\
        );

    \I__4198\ : InMux
    port map (
            O => \N__20789\,
            I => \N__20730\
        );

    \I__4197\ : InMux
    port map (
            O => \N__20786\,
            I => \N__20730\
        );

    \I__4196\ : InMux
    port map (
            O => \N__20783\,
            I => \N__20730\
        );

    \I__4195\ : InMux
    port map (
            O => \N__20780\,
            I => \N__20730\
        );

    \I__4194\ : InMux
    port map (
            O => \N__20777\,
            I => \N__20721\
        );

    \I__4193\ : InMux
    port map (
            O => \N__20774\,
            I => \N__20721\
        );

    \I__4192\ : InMux
    port map (
            O => \N__20771\,
            I => \N__20721\
        );

    \I__4191\ : InMux
    port map (
            O => \N__20768\,
            I => \N__20721\
        );

    \I__4190\ : InMux
    port map (
            O => \N__20767\,
            I => \N__20718\
        );

    \I__4189\ : LocalMux
    port map (
            O => \N__20764\,
            I => \N__20713\
        );

    \I__4188\ : Span4Mux_h
    port map (
            O => \N__20761\,
            I => \N__20713\
        );

    \I__4187\ : Span12Mux_s6_h
    port map (
            O => \N__20758\,
            I => \N__20710\
        );

    \I__4186\ : InMux
    port map (
            O => \N__20757\,
            I => \N__20705\
        );

    \I__4185\ : InMux
    port map (
            O => \N__20756\,
            I => \N__20705\
        );

    \I__4184\ : InMux
    port map (
            O => \N__20755\,
            I => \N__20698\
        );

    \I__4183\ : InMux
    port map (
            O => \N__20752\,
            I => \N__20698\
        );

    \I__4182\ : InMux
    port map (
            O => \N__20751\,
            I => \N__20698\
        );

    \I__4181\ : InMux
    port map (
            O => \N__20748\,
            I => \N__20685\
        );

    \I__4180\ : InMux
    port map (
            O => \N__20747\,
            I => \N__20685\
        );

    \I__4179\ : InMux
    port map (
            O => \N__20746\,
            I => \N__20685\
        );

    \I__4178\ : InMux
    port map (
            O => \N__20743\,
            I => \N__20685\
        );

    \I__4177\ : InMux
    port map (
            O => \N__20742\,
            I => \N__20685\
        );

    \I__4176\ : InMux
    port map (
            O => \N__20739\,
            I => \N__20685\
        );

    \I__4175\ : LocalMux
    port map (
            O => \N__20730\,
            I => \Lab_UT.dictrl.nextStateZ0Z_2\
        );

    \I__4174\ : LocalMux
    port map (
            O => \N__20721\,
            I => \Lab_UT.dictrl.nextStateZ0Z_2\
        );

    \I__4173\ : LocalMux
    port map (
            O => \N__20718\,
            I => \Lab_UT.dictrl.nextStateZ0Z_2\
        );

    \I__4172\ : Odrv4
    port map (
            O => \N__20713\,
            I => \Lab_UT.dictrl.nextStateZ0Z_2\
        );

    \I__4171\ : Odrv12
    port map (
            O => \N__20710\,
            I => \Lab_UT.dictrl.nextStateZ0Z_2\
        );

    \I__4170\ : LocalMux
    port map (
            O => \N__20705\,
            I => \Lab_UT.dictrl.nextStateZ0Z_2\
        );

    \I__4169\ : LocalMux
    port map (
            O => \N__20698\,
            I => \Lab_UT.dictrl.nextStateZ0Z_2\
        );

    \I__4168\ : LocalMux
    port map (
            O => \N__20685\,
            I => \Lab_UT.dictrl.nextStateZ0Z_2\
        );

    \I__4167\ : InMux
    port map (
            O => \N__20668\,
            I => \N__20654\
        );

    \I__4166\ : InMux
    port map (
            O => \N__20667\,
            I => \N__20644\
        );

    \I__4165\ : InMux
    port map (
            O => \N__20666\,
            I => \N__20644\
        );

    \I__4164\ : InMux
    port map (
            O => \N__20665\,
            I => \N__20644\
        );

    \I__4163\ : InMux
    port map (
            O => \N__20664\,
            I => \N__20644\
        );

    \I__4162\ : InMux
    port map (
            O => \N__20663\,
            I => \N__20635\
        );

    \I__4161\ : InMux
    port map (
            O => \N__20662\,
            I => \N__20635\
        );

    \I__4160\ : InMux
    port map (
            O => \N__20661\,
            I => \N__20635\
        );

    \I__4159\ : InMux
    port map (
            O => \N__20660\,
            I => \N__20635\
        );

    \I__4158\ : CascadeMux
    port map (
            O => \N__20659\,
            I => \N__20631\
        );

    \I__4157\ : CascadeMux
    port map (
            O => \N__20658\,
            I => \N__20628\
        );

    \I__4156\ : CascadeMux
    port map (
            O => \N__20657\,
            I => \N__20624\
        );

    \I__4155\ : LocalMux
    port map (
            O => \N__20654\,
            I => \N__20619\
        );

    \I__4154\ : InMux
    port map (
            O => \N__20653\,
            I => \N__20616\
        );

    \I__4153\ : LocalMux
    port map (
            O => \N__20644\,
            I => \N__20611\
        );

    \I__4152\ : LocalMux
    port map (
            O => \N__20635\,
            I => \N__20611\
        );

    \I__4151\ : InMux
    port map (
            O => \N__20634\,
            I => \N__20598\
        );

    \I__4150\ : InMux
    port map (
            O => \N__20631\,
            I => \N__20598\
        );

    \I__4149\ : InMux
    port map (
            O => \N__20628\,
            I => \N__20598\
        );

    \I__4148\ : InMux
    port map (
            O => \N__20627\,
            I => \N__20598\
        );

    \I__4147\ : InMux
    port map (
            O => \N__20624\,
            I => \N__20598\
        );

    \I__4146\ : InMux
    port map (
            O => \N__20623\,
            I => \N__20598\
        );

    \I__4145\ : InMux
    port map (
            O => \N__20622\,
            I => \N__20595\
        );

    \I__4144\ : Span4Mux_h
    port map (
            O => \N__20619\,
            I => \N__20592\
        );

    \I__4143\ : LocalMux
    port map (
            O => \N__20616\,
            I => \N__20585\
        );

    \I__4142\ : Span12Mux_s6_v
    port map (
            O => \N__20611\,
            I => \N__20585\
        );

    \I__4141\ : LocalMux
    port map (
            O => \N__20598\,
            I => \N__20585\
        );

    \I__4140\ : LocalMux
    port map (
            O => \N__20595\,
            I => \Lab_UT.dictrl.nextStateZ0Z_1\
        );

    \I__4139\ : Odrv4
    port map (
            O => \N__20592\,
            I => \Lab_UT.dictrl.nextStateZ0Z_1\
        );

    \I__4138\ : Odrv12
    port map (
            O => \N__20585\,
            I => \Lab_UT.dictrl.nextStateZ0Z_1\
        );

    \I__4137\ : InMux
    port map (
            O => \N__20578\,
            I => \N__20575\
        );

    \I__4136\ : LocalMux
    port map (
            O => \N__20575\,
            I => \N__20572\
        );

    \I__4135\ : Odrv4
    port map (
            O => \N__20572\,
            I => \Lab_UT.dictrl.r_dicLdMtens17\
        );

    \I__4134\ : InMux
    port map (
            O => \N__20569\,
            I => \N__20566\
        );

    \I__4133\ : LocalMux
    port map (
            O => \N__20566\,
            I => \N__20563\
        );

    \I__4132\ : Span4Mux_h
    port map (
            O => \N__20563\,
            I => \N__20557\
        );

    \I__4131\ : InMux
    port map (
            O => \N__20562\,
            I => \N__20554\
        );

    \I__4130\ : InMux
    port map (
            O => \N__20561\,
            I => \N__20551\
        );

    \I__4129\ : InMux
    port map (
            O => \N__20560\,
            I => \N__20548\
        );

    \I__4128\ : Odrv4
    port map (
            O => \N__20557\,
            I => \Lab_UT.dictrl.currState_ret_1and\
        );

    \I__4127\ : LocalMux
    port map (
            O => \N__20554\,
            I => \Lab_UT.dictrl.currState_ret_1and\
        );

    \I__4126\ : LocalMux
    port map (
            O => \N__20551\,
            I => \Lab_UT.dictrl.currState_ret_1and\
        );

    \I__4125\ : LocalMux
    port map (
            O => \N__20548\,
            I => \Lab_UT.dictrl.currState_ret_1and\
        );

    \I__4124\ : CascadeMux
    port map (
            O => \N__20539\,
            I => \N__20536\
        );

    \I__4123\ : InMux
    port map (
            O => \N__20536\,
            I => \N__20533\
        );

    \I__4122\ : LocalMux
    port map (
            O => \N__20533\,
            I => \Lab_UT.dictrl.dicLdAMones_rst\
        );

    \I__4121\ : InMux
    port map (
            O => \N__20530\,
            I => \N__20524\
        );

    \I__4120\ : InMux
    port map (
            O => \N__20529\,
            I => \N__20524\
        );

    \I__4119\ : LocalMux
    port map (
            O => \N__20524\,
            I => \Lab_UT.dictrl.dicLdAMonesZ0\
        );

    \I__4118\ : CascadeMux
    port map (
            O => \N__20521\,
            I => \Lab_UT.dictrl.dicLdAMones_rst_cascade_\
        );

    \I__4117\ : InMux
    port map (
            O => \N__20518\,
            I => \N__20508\
        );

    \I__4116\ : InMux
    port map (
            O => \N__20517\,
            I => \N__20508\
        );

    \I__4115\ : InMux
    port map (
            O => \N__20516\,
            I => \N__20508\
        );

    \I__4114\ : InMux
    port map (
            O => \N__20515\,
            I => \N__20503\
        );

    \I__4113\ : LocalMux
    port map (
            O => \N__20508\,
            I => \N__20500\
        );

    \I__4112\ : InMux
    port map (
            O => \N__20507\,
            I => \N__20495\
        );

    \I__4111\ : InMux
    port map (
            O => \N__20506\,
            I => \N__20495\
        );

    \I__4110\ : LocalMux
    port map (
            O => \N__20503\,
            I => \N__20492\
        );

    \I__4109\ : Span4Mux_h
    port map (
            O => \N__20500\,
            I => \N__20487\
        );

    \I__4108\ : LocalMux
    port map (
            O => \N__20495\,
            I => \N__20487\
        );

    \I__4107\ : Span4Mux_v
    port map (
            O => \N__20492\,
            I => \N__20484\
        );

    \I__4106\ : Span4Mux_v
    port map (
            O => \N__20487\,
            I => \N__20481\
        );

    \I__4105\ : Odrv4
    port map (
            O => \N__20484\,
            I => \Lab_UT.dictrl.r_dicLdMtens23_2\
        );

    \I__4104\ : Odrv4
    port map (
            O => \N__20481\,
            I => \Lab_UT.dictrl.r_dicLdMtens23_2\
        );

    \I__4103\ : CascadeMux
    port map (
            O => \N__20476\,
            I => \N__20472\
        );

    \I__4102\ : InMux
    port map (
            O => \N__20475\,
            I => \N__20469\
        );

    \I__4101\ : InMux
    port map (
            O => \N__20472\,
            I => \N__20466\
        );

    \I__4100\ : LocalMux
    port map (
            O => \N__20469\,
            I => \N__20463\
        );

    \I__4099\ : LocalMux
    port map (
            O => \N__20466\,
            I => \Lab_UT.dictrl.dicLdAStensZ0\
        );

    \I__4098\ : Odrv12
    port map (
            O => \N__20463\,
            I => \Lab_UT.dictrl.dicLdAStensZ0\
        );

    \I__4097\ : InMux
    port map (
            O => \N__20458\,
            I => \N__20454\
        );

    \I__4096\ : InMux
    port map (
            O => \N__20457\,
            I => \N__20451\
        );

    \I__4095\ : LocalMux
    port map (
            O => \N__20454\,
            I => \N__20448\
        );

    \I__4094\ : LocalMux
    port map (
            O => \N__20451\,
            I => \N__20445\
        );

    \I__4093\ : Span4Mux_v
    port map (
            O => \N__20448\,
            I => \N__20442\
        );

    \I__4092\ : Span4Mux_v
    port map (
            O => \N__20445\,
            I => \N__20437\
        );

    \I__4091\ : Span4Mux_h
    port map (
            O => \N__20442\,
            I => \N__20437\
        );

    \I__4090\ : Odrv4
    port map (
            O => \N__20437\,
            I => \Lab_UT.dictrl.dicLdAStens_rst\
        );

    \I__4089\ : InMux
    port map (
            O => \N__20434\,
            I => \N__20428\
        );

    \I__4088\ : InMux
    port map (
            O => \N__20433\,
            I => \N__20428\
        );

    \I__4087\ : LocalMux
    port map (
            O => \N__20428\,
            I => \N__20425\
        );

    \I__4086\ : Span4Mux_v
    port map (
            O => \N__20425\,
            I => \N__20419\
        );

    \I__4085\ : InMux
    port map (
            O => \N__20424\,
            I => \N__20412\
        );

    \I__4084\ : InMux
    port map (
            O => \N__20423\,
            I => \N__20412\
        );

    \I__4083\ : InMux
    port map (
            O => \N__20422\,
            I => \N__20412\
        );

    \I__4082\ : Sp12to4
    port map (
            O => \N__20419\,
            I => \N__20409\
        );

    \I__4081\ : LocalMux
    port map (
            O => \N__20412\,
            I => \N__20406\
        );

    \I__4080\ : Span12Mux_s7_h
    port map (
            O => \N__20409\,
            I => \N__20401\
        );

    \I__4079\ : Span12Mux_s4_v
    port map (
            O => \N__20406\,
            I => \N__20401\
        );

    \I__4078\ : Odrv12
    port map (
            O => \N__20401\,
            I => \resetGen.escKeyZ0\
        );

    \I__4077\ : CascadeMux
    port map (
            O => \N__20398\,
            I => \N__20389\
        );

    \I__4076\ : CascadeMux
    port map (
            O => \N__20397\,
            I => \N__20385\
        );

    \I__4075\ : CascadeMux
    port map (
            O => \N__20396\,
            I => \N__20382\
        );

    \I__4074\ : InMux
    port map (
            O => \N__20395\,
            I => \N__20379\
        );

    \I__4073\ : InMux
    port map (
            O => \N__20394\,
            I => \N__20374\
        );

    \I__4072\ : InMux
    port map (
            O => \N__20393\,
            I => \N__20374\
        );

    \I__4071\ : InMux
    port map (
            O => \N__20392\,
            I => \N__20371\
        );

    \I__4070\ : InMux
    port map (
            O => \N__20389\,
            I => \N__20362\
        );

    \I__4069\ : InMux
    port map (
            O => \N__20388\,
            I => \N__20362\
        );

    \I__4068\ : InMux
    port map (
            O => \N__20385\,
            I => \N__20362\
        );

    \I__4067\ : InMux
    port map (
            O => \N__20382\,
            I => \N__20357\
        );

    \I__4066\ : LocalMux
    port map (
            O => \N__20379\,
            I => \N__20352\
        );

    \I__4065\ : LocalMux
    port map (
            O => \N__20374\,
            I => \N__20352\
        );

    \I__4064\ : LocalMux
    port map (
            O => \N__20371\,
            I => \N__20349\
        );

    \I__4063\ : InMux
    port map (
            O => \N__20370\,
            I => \N__20346\
        );

    \I__4062\ : InMux
    port map (
            O => \N__20369\,
            I => \N__20343\
        );

    \I__4061\ : LocalMux
    port map (
            O => \N__20362\,
            I => \N__20340\
        );

    \I__4060\ : InMux
    port map (
            O => \N__20361\,
            I => \N__20335\
        );

    \I__4059\ : InMux
    port map (
            O => \N__20360\,
            I => \N__20335\
        );

    \I__4058\ : LocalMux
    port map (
            O => \N__20357\,
            I => \N__20329\
        );

    \I__4057\ : Span4Mux_v
    port map (
            O => \N__20352\,
            I => \N__20329\
        );

    \I__4056\ : Span4Mux_v
    port map (
            O => \N__20349\,
            I => \N__20324\
        );

    \I__4055\ : LocalMux
    port map (
            O => \N__20346\,
            I => \N__20324\
        );

    \I__4054\ : LocalMux
    port map (
            O => \N__20343\,
            I => \N__20321\
        );

    \I__4053\ : Span4Mux_h
    port map (
            O => \N__20340\,
            I => \N__20316\
        );

    \I__4052\ : LocalMux
    port map (
            O => \N__20335\,
            I => \N__20316\
        );

    \I__4051\ : InMux
    port map (
            O => \N__20334\,
            I => \N__20313\
        );

    \I__4050\ : Span4Mux_h
    port map (
            O => \N__20329\,
            I => \N__20308\
        );

    \I__4049\ : Span4Mux_v
    port map (
            O => \N__20324\,
            I => \N__20308\
        );

    \I__4048\ : Odrv4
    port map (
            O => \N__20321\,
            I => \Lab_UT.dictrl.currState_3_rep1\
        );

    \I__4047\ : Odrv4
    port map (
            O => \N__20316\,
            I => \Lab_UT.dictrl.currState_3_rep1\
        );

    \I__4046\ : LocalMux
    port map (
            O => \N__20313\,
            I => \Lab_UT.dictrl.currState_3_rep1\
        );

    \I__4045\ : Odrv4
    port map (
            O => \N__20308\,
            I => \Lab_UT.dictrl.currState_3_rep1\
        );

    \I__4044\ : InMux
    port map (
            O => \N__20299\,
            I => \N__20296\
        );

    \I__4043\ : LocalMux
    port map (
            O => \N__20296\,
            I => \N__20292\
        );

    \I__4042\ : InMux
    port map (
            O => \N__20295\,
            I => \N__20289\
        );

    \I__4041\ : Odrv12
    port map (
            O => \N__20292\,
            I => \Lab_UT.dictrl.N_5\
        );

    \I__4040\ : LocalMux
    port map (
            O => \N__20289\,
            I => \Lab_UT.dictrl.N_5\
        );

    \I__4039\ : InMux
    port map (
            O => \N__20284\,
            I => \N__20280\
        );

    \I__4038\ : InMux
    port map (
            O => \N__20283\,
            I => \N__20277\
        );

    \I__4037\ : LocalMux
    port map (
            O => \N__20280\,
            I => \N__20274\
        );

    \I__4036\ : LocalMux
    port map (
            O => \N__20277\,
            I => \N__20271\
        );

    \I__4035\ : Span4Mux_h
    port map (
            O => \N__20274\,
            I => \N__20268\
        );

    \I__4034\ : Odrv4
    port map (
            O => \N__20271\,
            I => \Lab_UT.dictrl.N_6\
        );

    \I__4033\ : Odrv4
    port map (
            O => \N__20268\,
            I => \Lab_UT.dictrl.N_6\
        );

    \I__4032\ : CascadeMux
    port map (
            O => \N__20263\,
            I => \Lab_UT.dictrl.r_enable2_3_iv_0_cascade_\
        );

    \I__4031\ : InMux
    port map (
            O => \N__20260\,
            I => \N__20257\
        );

    \I__4030\ : LocalMux
    port map (
            O => \N__20257\,
            I => \N__20254\
        );

    \I__4029\ : Odrv4
    port map (
            O => \N__20254\,
            I => \Lab_UT.dictrl.r_enable2_3_iv_3\
        );

    \I__4028\ : InMux
    port map (
            O => \N__20251\,
            I => \N__20248\
        );

    \I__4027\ : LocalMux
    port map (
            O => \N__20248\,
            I => \N__20245\
        );

    \I__4026\ : Span4Mux_h
    port map (
            O => \N__20245\,
            I => \N__20242\
        );

    \I__4025\ : Sp12to4
    port map (
            O => \N__20242\,
            I => \N__20239\
        );

    \I__4024\ : Odrv12
    port map (
            O => \N__20239\,
            I => \Lab_UT.dictrl.r_Sone_init17_4\
        );

    \I__4023\ : InMux
    port map (
            O => \N__20236\,
            I => \N__20230\
        );

    \I__4022\ : InMux
    port map (
            O => \N__20235\,
            I => \N__20230\
        );

    \I__4021\ : LocalMux
    port map (
            O => \N__20230\,
            I => \Lab_UT.dictrl.r_dicLdMtens23_i_6\
        );

    \I__4020\ : CascadeMux
    port map (
            O => \N__20227\,
            I => \Lab_UT.dictrl.un1_r_dicLdMtens19_0_cascade_\
        );

    \I__4019\ : InMux
    port map (
            O => \N__20224\,
            I => \N__20220\
        );

    \I__4018\ : InMux
    port map (
            O => \N__20223\,
            I => \N__20217\
        );

    \I__4017\ : LocalMux
    port map (
            O => \N__20220\,
            I => \Lab_UT.dictrl.r_alarm_or_timeZ0\
        );

    \I__4016\ : LocalMux
    port map (
            O => \N__20217\,
            I => \Lab_UT.dictrl.r_alarm_or_timeZ0\
        );

    \I__4015\ : InMux
    port map (
            O => \N__20212\,
            I => \N__20209\
        );

    \I__4014\ : LocalMux
    port map (
            O => \N__20209\,
            I => \Lab_UT.dictrl.r_dicLdMtens18_i_6\
        );

    \I__4013\ : InMux
    port map (
            O => \N__20206\,
            I => \N__20203\
        );

    \I__4012\ : LocalMux
    port map (
            O => \N__20203\,
            I => \Lab_UT.dictrl.r_dicLdMtens17_i_6\
        );

    \I__4011\ : InMux
    port map (
            O => \N__20200\,
            I => \N__20197\
        );

    \I__4010\ : LocalMux
    port map (
            O => \N__20197\,
            I => \N__20194\
        );

    \I__4009\ : Odrv4
    port map (
            O => \N__20194\,
            I => \Lab_UT.dictrl.r_enable1_2_m\
        );

    \I__4008\ : CascadeMux
    port map (
            O => \N__20191\,
            I => \Lab_UT.dictrl.r_enable1_2_m_cascade_\
        );

    \I__4007\ : InMux
    port map (
            O => \N__20188\,
            I => \N__20185\
        );

    \I__4006\ : LocalMux
    port map (
            O => \N__20185\,
            I => \N__20182\
        );

    \I__4005\ : Odrv12
    port map (
            O => \N__20182\,
            I => \Lab_UT.dictrl.g0_i_a4_0\
        );

    \I__4004\ : InMux
    port map (
            O => \N__20179\,
            I => \N__20173\
        );

    \I__4003\ : InMux
    port map (
            O => \N__20178\,
            I => \N__20173\
        );

    \I__4002\ : LocalMux
    port map (
            O => \N__20173\,
            I => \Lab_UT.dictrl.r_enableZ0Z2\
        );

    \I__4001\ : InMux
    port map (
            O => \N__20170\,
            I => \N__20161\
        );

    \I__4000\ : InMux
    port map (
            O => \N__20169\,
            I => \N__20154\
        );

    \I__3999\ : InMux
    port map (
            O => \N__20168\,
            I => \N__20154\
        );

    \I__3998\ : InMux
    port map (
            O => \N__20167\,
            I => \N__20154\
        );

    \I__3997\ : InMux
    port map (
            O => \N__20166\,
            I => \N__20147\
        );

    \I__3996\ : InMux
    port map (
            O => \N__20165\,
            I => \N__20147\
        );

    \I__3995\ : InMux
    port map (
            O => \N__20164\,
            I => \N__20147\
        );

    \I__3994\ : LocalMux
    port map (
            O => \N__20161\,
            I => \N__20144\
        );

    \I__3993\ : LocalMux
    port map (
            O => \N__20154\,
            I => \N__20141\
        );

    \I__3992\ : LocalMux
    port map (
            O => \N__20147\,
            I => \N__20138\
        );

    \I__3991\ : Span4Mux_v
    port map (
            O => \N__20144\,
            I => \N__20135\
        );

    \I__3990\ : Span4Mux_v
    port map (
            O => \N__20141\,
            I => \N__20130\
        );

    \I__3989\ : Span4Mux_h
    port map (
            O => \N__20138\,
            I => \N__20130\
        );

    \I__3988\ : Odrv4
    port map (
            O => \N__20135\,
            I => \Lab_UT.dictrl.enableSeg2\
        );

    \I__3987\ : Odrv4
    port map (
            O => \N__20130\,
            I => \Lab_UT.dictrl.enableSeg2\
        );

    \I__3986\ : InMux
    port map (
            O => \N__20125\,
            I => \N__20122\
        );

    \I__3985\ : LocalMux
    port map (
            O => \N__20122\,
            I => \Lab_UT.dictrl.currState_0_ret_20and_1_0\
        );

    \I__3984\ : InMux
    port map (
            O => \N__20119\,
            I => \N__20115\
        );

    \I__3983\ : InMux
    port map (
            O => \N__20118\,
            I => \N__20112\
        );

    \I__3982\ : LocalMux
    port map (
            O => \N__20115\,
            I => \Lab_UT.dictrl.r_dicLdMtens16_reti\
        );

    \I__3981\ : LocalMux
    port map (
            O => \N__20112\,
            I => \Lab_UT.dictrl.r_dicLdMtens16_reti\
        );

    \I__3980\ : InMux
    port map (
            O => \N__20107\,
            I => \N__20103\
        );

    \I__3979\ : InMux
    port map (
            O => \N__20106\,
            I => \N__20100\
        );

    \I__3978\ : LocalMux
    port map (
            O => \N__20103\,
            I => \N__20095\
        );

    \I__3977\ : LocalMux
    port map (
            O => \N__20100\,
            I => \N__20095\
        );

    \I__3976\ : Span4Mux_v
    port map (
            O => \N__20095\,
            I => \N__20092\
        );

    \I__3975\ : Span4Mux_h
    port map (
            O => \N__20092\,
            I => \N__20089\
        );

    \I__3974\ : Odrv4
    port map (
            O => \N__20089\,
            I => \Lab_UT.dictrl.r_dicLdMtens19\
        );

    \I__3973\ : InMux
    port map (
            O => \N__20086\,
            I => \N__20083\
        );

    \I__3972\ : LocalMux
    port map (
            O => \N__20083\,
            I => \N__20080\
        );

    \I__3971\ : Odrv12
    port map (
            O => \N__20080\,
            I => \Lab_UT.dictrl.r_dicLdMtens22_i_6\
        );

    \I__3970\ : InMux
    port map (
            O => \N__20077\,
            I => \N__20062\
        );

    \I__3969\ : InMux
    port map (
            O => \N__20076\,
            I => \N__20062\
        );

    \I__3968\ : InMux
    port map (
            O => \N__20075\,
            I => \N__20062\
        );

    \I__3967\ : InMux
    port map (
            O => \N__20074\,
            I => \N__20062\
        );

    \I__3966\ : InMux
    port map (
            O => \N__20073\,
            I => \N__20055\
        );

    \I__3965\ : InMux
    port map (
            O => \N__20072\,
            I => \N__20055\
        );

    \I__3964\ : InMux
    port map (
            O => \N__20071\,
            I => \N__20055\
        );

    \I__3963\ : LocalMux
    port map (
            O => \N__20062\,
            I => \N__20052\
        );

    \I__3962\ : LocalMux
    port map (
            O => \N__20055\,
            I => \Lab_UT.Sten_at_1\
        );

    \I__3961\ : Odrv4
    port map (
            O => \N__20052\,
            I => \Lab_UT.Sten_at_1\
        );

    \I__3960\ : InMux
    port map (
            O => \N__20047\,
            I => \N__20031\
        );

    \I__3959\ : InMux
    port map (
            O => \N__20046\,
            I => \N__20031\
        );

    \I__3958\ : InMux
    port map (
            O => \N__20045\,
            I => \N__20031\
        );

    \I__3957\ : InMux
    port map (
            O => \N__20044\,
            I => \N__20031\
        );

    \I__3956\ : InMux
    port map (
            O => \N__20043\,
            I => \N__20021\
        );

    \I__3955\ : InMux
    port map (
            O => \N__20042\,
            I => \N__20021\
        );

    \I__3954\ : InMux
    port map (
            O => \N__20041\,
            I => \N__20021\
        );

    \I__3953\ : InMux
    port map (
            O => \N__20040\,
            I => \N__20021\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__20031\,
            I => \N__20018\
        );

    \I__3951\ : InMux
    port map (
            O => \N__20030\,
            I => \N__20015\
        );

    \I__3950\ : LocalMux
    port map (
            O => \N__20021\,
            I => \Lab_UT.Sten_at_0\
        );

    \I__3949\ : Odrv4
    port map (
            O => \N__20018\,
            I => \Lab_UT.Sten_at_0\
        );

    \I__3948\ : LocalMux
    port map (
            O => \N__20015\,
            I => \Lab_UT.Sten_at_0\
        );

    \I__3947\ : CascadeMux
    port map (
            O => \N__20008\,
            I => \N__20002\
        );

    \I__3946\ : InMux
    port map (
            O => \N__20007\,
            I => \N__19993\
        );

    \I__3945\ : InMux
    port map (
            O => \N__20006\,
            I => \N__19993\
        );

    \I__3944\ : InMux
    port map (
            O => \N__20005\,
            I => \N__19993\
        );

    \I__3943\ : InMux
    port map (
            O => \N__20002\,
            I => \N__19993\
        );

    \I__3942\ : LocalMux
    port map (
            O => \N__19993\,
            I => \N__19988\
        );

    \I__3941\ : CascadeMux
    port map (
            O => \N__19992\,
            I => \N__19984\
        );

    \I__3940\ : CascadeMux
    port map (
            O => \N__19991\,
            I => \N__19980\
        );

    \I__3939\ : Span4Mux_h
    port map (
            O => \N__19988\,
            I => \N__19976\
        );

    \I__3938\ : InMux
    port map (
            O => \N__19987\,
            I => \N__19973\
        );

    \I__3937\ : InMux
    port map (
            O => \N__19984\,
            I => \N__19966\
        );

    \I__3936\ : InMux
    port map (
            O => \N__19983\,
            I => \N__19966\
        );

    \I__3935\ : InMux
    port map (
            O => \N__19980\,
            I => \N__19966\
        );

    \I__3934\ : InMux
    port map (
            O => \N__19979\,
            I => \N__19963\
        );

    \I__3933\ : Odrv4
    port map (
            O => \N__19976\,
            I => \Lab_UT.Sten_at_3\
        );

    \I__3932\ : LocalMux
    port map (
            O => \N__19973\,
            I => \Lab_UT.Sten_at_3\
        );

    \I__3931\ : LocalMux
    port map (
            O => \N__19966\,
            I => \Lab_UT.Sten_at_3\
        );

    \I__3930\ : LocalMux
    port map (
            O => \N__19963\,
            I => \Lab_UT.Sten_at_3\
        );

    \I__3929\ : CascadeMux
    port map (
            O => \N__19954\,
            I => \Lab_UT.Sten_at_1_cascade_\
        );

    \I__3928\ : CascadeMux
    port map (
            O => \N__19951\,
            I => \N__19945\
        );

    \I__3927\ : CascadeMux
    port map (
            O => \N__19950\,
            I => \N__19942\
        );

    \I__3926\ : CascadeMux
    port map (
            O => \N__19949\,
            I => \N__19939\
        );

    \I__3925\ : CascadeMux
    port map (
            O => \N__19948\,
            I => \N__19934\
        );

    \I__3924\ : InMux
    port map (
            O => \N__19945\,
            I => \N__19924\
        );

    \I__3923\ : InMux
    port map (
            O => \N__19942\,
            I => \N__19924\
        );

    \I__3922\ : InMux
    port map (
            O => \N__19939\,
            I => \N__19924\
        );

    \I__3921\ : InMux
    port map (
            O => \N__19938\,
            I => \N__19924\
        );

    \I__3920\ : InMux
    port map (
            O => \N__19937\,
            I => \N__19916\
        );

    \I__3919\ : InMux
    port map (
            O => \N__19934\,
            I => \N__19916\
        );

    \I__3918\ : InMux
    port map (
            O => \N__19933\,
            I => \N__19916\
        );

    \I__3917\ : LocalMux
    port map (
            O => \N__19924\,
            I => \N__19913\
        );

    \I__3916\ : InMux
    port map (
            O => \N__19923\,
            I => \N__19910\
        );

    \I__3915\ : LocalMux
    port map (
            O => \N__19916\,
            I => \Lab_UT.Sten_at_2\
        );

    \I__3914\ : Odrv4
    port map (
            O => \N__19913\,
            I => \Lab_UT.Sten_at_2\
        );

    \I__3913\ : LocalMux
    port map (
            O => \N__19910\,
            I => \Lab_UT.Sten_at_2\
        );

    \I__3912\ : InMux
    port map (
            O => \N__19903\,
            I => \N__19900\
        );

    \I__3911\ : LocalMux
    port map (
            O => \N__19900\,
            I => \Lab_UT.segmentUQ_0_0_0\
        );

    \I__3910\ : CascadeMux
    port map (
            O => \N__19897\,
            I => \N__19890\
        );

    \I__3909\ : InMux
    port map (
            O => \N__19896\,
            I => \N__19870\
        );

    \I__3908\ : InMux
    port map (
            O => \N__19895\,
            I => \N__19870\
        );

    \I__3907\ : InMux
    port map (
            O => \N__19894\,
            I => \N__19865\
        );

    \I__3906\ : InMux
    port map (
            O => \N__19893\,
            I => \N__19865\
        );

    \I__3905\ : InMux
    port map (
            O => \N__19890\,
            I => \N__19858\
        );

    \I__3904\ : InMux
    port map (
            O => \N__19889\,
            I => \N__19858\
        );

    \I__3903\ : InMux
    port map (
            O => \N__19888\,
            I => \N__19858\
        );

    \I__3902\ : CascadeMux
    port map (
            O => \N__19887\,
            I => \N__19852\
        );

    \I__3901\ : InMux
    port map (
            O => \N__19886\,
            I => \N__19845\
        );

    \I__3900\ : InMux
    port map (
            O => \N__19885\,
            I => \N__19840\
        );

    \I__3899\ : InMux
    port map (
            O => \N__19884\,
            I => \N__19840\
        );

    \I__3898\ : InMux
    port map (
            O => \N__19883\,
            I => \N__19835\
        );

    \I__3897\ : InMux
    port map (
            O => \N__19882\,
            I => \N__19835\
        );

    \I__3896\ : InMux
    port map (
            O => \N__19881\,
            I => \N__19828\
        );

    \I__3895\ : InMux
    port map (
            O => \N__19880\,
            I => \N__19828\
        );

    \I__3894\ : InMux
    port map (
            O => \N__19879\,
            I => \N__19828\
        );

    \I__3893\ : InMux
    port map (
            O => \N__19878\,
            I => \N__19821\
        );

    \I__3892\ : InMux
    port map (
            O => \N__19877\,
            I => \N__19821\
        );

    \I__3891\ : InMux
    port map (
            O => \N__19876\,
            I => \N__19821\
        );

    \I__3890\ : CascadeMux
    port map (
            O => \N__19875\,
            I => \N__19817\
        );

    \I__3889\ : LocalMux
    port map (
            O => \N__19870\,
            I => \N__19810\
        );

    \I__3888\ : LocalMux
    port map (
            O => \N__19865\,
            I => \N__19810\
        );

    \I__3887\ : LocalMux
    port map (
            O => \N__19858\,
            I => \N__19810\
        );

    \I__3886\ : InMux
    port map (
            O => \N__19857\,
            I => \N__19807\
        );

    \I__3885\ : InMux
    port map (
            O => \N__19856\,
            I => \N__19802\
        );

    \I__3884\ : InMux
    port map (
            O => \N__19855\,
            I => \N__19802\
        );

    \I__3883\ : InMux
    port map (
            O => \N__19852\,
            I => \N__19797\
        );

    \I__3882\ : InMux
    port map (
            O => \N__19851\,
            I => \N__19797\
        );

    \I__3881\ : InMux
    port map (
            O => \N__19850\,
            I => \N__19790\
        );

    \I__3880\ : InMux
    port map (
            O => \N__19849\,
            I => \N__19790\
        );

    \I__3879\ : InMux
    port map (
            O => \N__19848\,
            I => \N__19790\
        );

    \I__3878\ : LocalMux
    port map (
            O => \N__19845\,
            I => \N__19783\
        );

    \I__3877\ : LocalMux
    port map (
            O => \N__19840\,
            I => \N__19783\
        );

    \I__3876\ : LocalMux
    port map (
            O => \N__19835\,
            I => \N__19783\
        );

    \I__3875\ : LocalMux
    port map (
            O => \N__19828\,
            I => \N__19778\
        );

    \I__3874\ : LocalMux
    port map (
            O => \N__19821\,
            I => \N__19778\
        );

    \I__3873\ : InMux
    port map (
            O => \N__19820\,
            I => \N__19773\
        );

    \I__3872\ : InMux
    port map (
            O => \N__19817\,
            I => \N__19773\
        );

    \I__3871\ : Span4Mux_v
    port map (
            O => \N__19810\,
            I => \N__19770\
        );

    \I__3870\ : LocalMux
    port map (
            O => \N__19807\,
            I => \N__19761\
        );

    \I__3869\ : LocalMux
    port map (
            O => \N__19802\,
            I => \N__19761\
        );

    \I__3868\ : LocalMux
    port map (
            O => \N__19797\,
            I => \N__19761\
        );

    \I__3867\ : LocalMux
    port map (
            O => \N__19790\,
            I => \N__19761\
        );

    \I__3866\ : Span4Mux_h
    port map (
            O => \N__19783\,
            I => \N__19758\
        );

    \I__3865\ : Span4Mux_h
    port map (
            O => \N__19778\,
            I => \N__19755\
        );

    \I__3864\ : LocalMux
    port map (
            O => \N__19773\,
            I => \N__19750\
        );

    \I__3863\ : Span4Mux_h
    port map (
            O => \N__19770\,
            I => \N__19750\
        );

    \I__3862\ : Odrv4
    port map (
            O => \N__19761\,
            I => \Lab_UT.dictrl.L3_segment1_1\
        );

    \I__3861\ : Odrv4
    port map (
            O => \N__19758\,
            I => \Lab_UT.dictrl.L3_segment1_1\
        );

    \I__3860\ : Odrv4
    port map (
            O => \N__19755\,
            I => \Lab_UT.dictrl.L3_segment1_1\
        );

    \I__3859\ : Odrv4
    port map (
            O => \N__19750\,
            I => \Lab_UT.dictrl.L3_segment1_1\
        );

    \I__3858\ : CascadeMux
    port map (
            O => \N__19741\,
            I => \N__19733\
        );

    \I__3857\ : CascadeMux
    port map (
            O => \N__19740\,
            I => \N__19730\
        );

    \I__3856\ : CascadeMux
    port map (
            O => \N__19739\,
            I => \N__19727\
        );

    \I__3855\ : CascadeMux
    port map (
            O => \N__19738\,
            I => \N__19723\
        );

    \I__3854\ : InMux
    port map (
            O => \N__19737\,
            I => \N__19713\
        );

    \I__3853\ : InMux
    port map (
            O => \N__19736\,
            I => \N__19713\
        );

    \I__3852\ : InMux
    port map (
            O => \N__19733\,
            I => \N__19713\
        );

    \I__3851\ : InMux
    port map (
            O => \N__19730\,
            I => \N__19713\
        );

    \I__3850\ : InMux
    port map (
            O => \N__19727\,
            I => \N__19704\
        );

    \I__3849\ : InMux
    port map (
            O => \N__19726\,
            I => \N__19704\
        );

    \I__3848\ : InMux
    port map (
            O => \N__19723\,
            I => \N__19704\
        );

    \I__3847\ : InMux
    port map (
            O => \N__19722\,
            I => \N__19704\
        );

    \I__3846\ : LocalMux
    port map (
            O => \N__19713\,
            I => \N__19699\
        );

    \I__3845\ : LocalMux
    port map (
            O => \N__19704\,
            I => \N__19699\
        );

    \I__3844\ : Odrv4
    port map (
            O => \N__19699\,
            I => \Lab_UT.Sone_at_1\
        );

    \I__3843\ : InMux
    port map (
            O => \N__19696\,
            I => \N__19690\
        );

    \I__3842\ : InMux
    port map (
            O => \N__19695\,
            I => \N__19690\
        );

    \I__3841\ : LocalMux
    port map (
            O => \N__19690\,
            I => \N__19687\
        );

    \I__3840\ : Odrv4
    port map (
            O => \N__19687\,
            I => \Lab_UT.dictrl.r_enable1_2_i_m\
        );

    \I__3839\ : InMux
    port map (
            O => \N__19684\,
            I => \N__19672\
        );

    \I__3838\ : InMux
    port map (
            O => \N__19683\,
            I => \N__19672\
        );

    \I__3837\ : InMux
    port map (
            O => \N__19682\,
            I => \N__19672\
        );

    \I__3836\ : InMux
    port map (
            O => \N__19681\,
            I => \N__19672\
        );

    \I__3835\ : LocalMux
    port map (
            O => \N__19672\,
            I => \N__19661\
        );

    \I__3834\ : InMux
    port map (
            O => \N__19671\,
            I => \N__19646\
        );

    \I__3833\ : InMux
    port map (
            O => \N__19670\,
            I => \N__19646\
        );

    \I__3832\ : InMux
    port map (
            O => \N__19669\,
            I => \N__19646\
        );

    \I__3831\ : InMux
    port map (
            O => \N__19668\,
            I => \N__19646\
        );

    \I__3830\ : InMux
    port map (
            O => \N__19667\,
            I => \N__19646\
        );

    \I__3829\ : InMux
    port map (
            O => \N__19666\,
            I => \N__19646\
        );

    \I__3828\ : InMux
    port map (
            O => \N__19665\,
            I => \N__19639\
        );

    \I__3827\ : InMux
    port map (
            O => \N__19664\,
            I => \N__19639\
        );

    \I__3826\ : Span4Mux_v
    port map (
            O => \N__19661\,
            I => \N__19636\
        );

    \I__3825\ : InMux
    port map (
            O => \N__19660\,
            I => \N__19631\
        );

    \I__3824\ : InMux
    port map (
            O => \N__19659\,
            I => \N__19631\
        );

    \I__3823\ : LocalMux
    port map (
            O => \N__19646\,
            I => \N__19628\
        );

    \I__3822\ : InMux
    port map (
            O => \N__19645\,
            I => \N__19623\
        );

    \I__3821\ : InMux
    port map (
            O => \N__19644\,
            I => \N__19623\
        );

    \I__3820\ : LocalMux
    port map (
            O => \N__19639\,
            I => \Lab_UT.alarm_or_time_0\
        );

    \I__3819\ : Odrv4
    port map (
            O => \N__19636\,
            I => \Lab_UT.alarm_or_time_0\
        );

    \I__3818\ : LocalMux
    port map (
            O => \N__19631\,
            I => \Lab_UT.alarm_or_time_0\
        );

    \I__3817\ : Odrv4
    port map (
            O => \N__19628\,
            I => \Lab_UT.alarm_or_time_0\
        );

    \I__3816\ : LocalMux
    port map (
            O => \N__19623\,
            I => \Lab_UT.alarm_or_time_0\
        );

    \I__3815\ : CascadeMux
    port map (
            O => \N__19612\,
            I => \Lab_UT.alarm_or_time_0_cascade_\
        );

    \I__3814\ : CascadeMux
    port map (
            O => \N__19609\,
            I => \N__19605\
        );

    \I__3813\ : InMux
    port map (
            O => \N__19608\,
            I => \N__19594\
        );

    \I__3812\ : InMux
    port map (
            O => \N__19605\,
            I => \N__19594\
        );

    \I__3811\ : InMux
    port map (
            O => \N__19604\,
            I => \N__19594\
        );

    \I__3810\ : InMux
    port map (
            O => \N__19603\,
            I => \N__19594\
        );

    \I__3809\ : LocalMux
    port map (
            O => \N__19594\,
            I => \N__19591\
        );

    \I__3808\ : Span4Mux_h
    port map (
            O => \N__19591\,
            I => \N__19584\
        );

    \I__3807\ : InMux
    port map (
            O => \N__19590\,
            I => \N__19581\
        );

    \I__3806\ : InMux
    port map (
            O => \N__19589\,
            I => \N__19576\
        );

    \I__3805\ : InMux
    port map (
            O => \N__19588\,
            I => \N__19576\
        );

    \I__3804\ : InMux
    port map (
            O => \N__19587\,
            I => \N__19573\
        );

    \I__3803\ : Odrv4
    port map (
            O => \N__19584\,
            I => \Lab_UT.Mten_at_2\
        );

    \I__3802\ : LocalMux
    port map (
            O => \N__19581\,
            I => \Lab_UT.Mten_at_2\
        );

    \I__3801\ : LocalMux
    port map (
            O => \N__19576\,
            I => \Lab_UT.Mten_at_2\
        );

    \I__3800\ : LocalMux
    port map (
            O => \N__19573\,
            I => \Lab_UT.Mten_at_2\
        );

    \I__3799\ : InMux
    port map (
            O => \N__19564\,
            I => \N__19556\
        );

    \I__3798\ : InMux
    port map (
            O => \N__19563\,
            I => \N__19549\
        );

    \I__3797\ : InMux
    port map (
            O => \N__19562\,
            I => \N__19549\
        );

    \I__3796\ : InMux
    port map (
            O => \N__19561\,
            I => \N__19549\
        );

    \I__3795\ : InMux
    port map (
            O => \N__19560\,
            I => \N__19544\
        );

    \I__3794\ : InMux
    port map (
            O => \N__19559\,
            I => \N__19544\
        );

    \I__3793\ : LocalMux
    port map (
            O => \N__19556\,
            I => \N__19536\
        );

    \I__3792\ : LocalMux
    port map (
            O => \N__19549\,
            I => \N__19536\
        );

    \I__3791\ : LocalMux
    port map (
            O => \N__19544\,
            I => \N__19536\
        );

    \I__3790\ : InMux
    port map (
            O => \N__19543\,
            I => \N__19533\
        );

    \I__3789\ : Span4Mux_h
    port map (
            O => \N__19536\,
            I => \N__19530\
        );

    \I__3788\ : LocalMux
    port map (
            O => \N__19533\,
            I => \N__19527\
        );

    \I__3787\ : Odrv4
    port map (
            O => \N__19530\,
            I => \Lab_UT.dictrl.enableSeg1\
        );

    \I__3786\ : Odrv12
    port map (
            O => \N__19527\,
            I => \Lab_UT.dictrl.enableSeg1\
        );

    \I__3785\ : CascadeMux
    port map (
            O => \N__19522\,
            I => \Lab_UT.L3_segment1_1_2_cascade_\
        );

    \I__3784\ : InMux
    port map (
            O => \N__19519\,
            I => \N__19516\
        );

    \I__3783\ : LocalMux
    port map (
            O => \N__19516\,
            I => \uu2.bitmapZ0Z_93\
        );

    \I__3782\ : InMux
    port map (
            O => \N__19513\,
            I => \N__19510\
        );

    \I__3781\ : LocalMux
    port map (
            O => \N__19510\,
            I => \uu2.bitmap_pmux_25_bm_1\
        );

    \I__3780\ : CascadeMux
    port map (
            O => \N__19507\,
            I => \N__19504\
        );

    \I__3779\ : InMux
    port map (
            O => \N__19504\,
            I => \N__19501\
        );

    \I__3778\ : LocalMux
    port map (
            O => \N__19501\,
            I => \uu2.bitmapZ0Z_221\
        );

    \I__3777\ : CascadeMux
    port map (
            O => \N__19498\,
            I => \N__19488\
        );

    \I__3776\ : CascadeMux
    port map (
            O => \N__19497\,
            I => \N__19484\
        );

    \I__3775\ : InMux
    port map (
            O => \N__19496\,
            I => \N__19480\
        );

    \I__3774\ : InMux
    port map (
            O => \N__19495\,
            I => \N__19477\
        );

    \I__3773\ : InMux
    port map (
            O => \N__19494\,
            I => \N__19474\
        );

    \I__3772\ : InMux
    port map (
            O => \N__19493\,
            I => \N__19468\
        );

    \I__3771\ : InMux
    port map (
            O => \N__19492\,
            I => \N__19468\
        );

    \I__3770\ : InMux
    port map (
            O => \N__19491\,
            I => \N__19465\
        );

    \I__3769\ : InMux
    port map (
            O => \N__19488\,
            I => \N__19460\
        );

    \I__3768\ : InMux
    port map (
            O => \N__19487\,
            I => \N__19460\
        );

    \I__3767\ : InMux
    port map (
            O => \N__19484\,
            I => \N__19453\
        );

    \I__3766\ : InMux
    port map (
            O => \N__19483\,
            I => \N__19453\
        );

    \I__3765\ : LocalMux
    port map (
            O => \N__19480\,
            I => \N__19448\
        );

    \I__3764\ : LocalMux
    port map (
            O => \N__19477\,
            I => \N__19448\
        );

    \I__3763\ : LocalMux
    port map (
            O => \N__19474\,
            I => \N__19445\
        );

    \I__3762\ : InMux
    port map (
            O => \N__19473\,
            I => \N__19442\
        );

    \I__3761\ : LocalMux
    port map (
            O => \N__19468\,
            I => \N__19439\
        );

    \I__3760\ : LocalMux
    port map (
            O => \N__19465\,
            I => \N__19432\
        );

    \I__3759\ : LocalMux
    port map (
            O => \N__19460\,
            I => \N__19429\
        );

    \I__3758\ : CascadeMux
    port map (
            O => \N__19459\,
            I => \N__19426\
        );

    \I__3757\ : CascadeMux
    port map (
            O => \N__19458\,
            I => \N__19422\
        );

    \I__3756\ : LocalMux
    port map (
            O => \N__19453\,
            I => \N__19415\
        );

    \I__3755\ : Span4Mux_h
    port map (
            O => \N__19448\,
            I => \N__19415\
        );

    \I__3754\ : Span4Mux_h
    port map (
            O => \N__19445\,
            I => \N__19415\
        );

    \I__3753\ : LocalMux
    port map (
            O => \N__19442\,
            I => \N__19410\
        );

    \I__3752\ : Span4Mux_h
    port map (
            O => \N__19439\,
            I => \N__19410\
        );

    \I__3751\ : InMux
    port map (
            O => \N__19438\,
            I => \N__19407\
        );

    \I__3750\ : InMux
    port map (
            O => \N__19437\,
            I => \N__19402\
        );

    \I__3749\ : InMux
    port map (
            O => \N__19436\,
            I => \N__19402\
        );

    \I__3748\ : InMux
    port map (
            O => \N__19435\,
            I => \N__19399\
        );

    \I__3747\ : Span4Mux_h
    port map (
            O => \N__19432\,
            I => \N__19394\
        );

    \I__3746\ : Span4Mux_h
    port map (
            O => \N__19429\,
            I => \N__19394\
        );

    \I__3745\ : InMux
    port map (
            O => \N__19426\,
            I => \N__19391\
        );

    \I__3744\ : InMux
    port map (
            O => \N__19425\,
            I => \N__19386\
        );

    \I__3743\ : InMux
    port map (
            O => \N__19422\,
            I => \N__19386\
        );

    \I__3742\ : Odrv4
    port map (
            O => \N__19415\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__3741\ : Odrv4
    port map (
            O => \N__19410\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__3740\ : LocalMux
    port map (
            O => \N__19407\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__3739\ : LocalMux
    port map (
            O => \N__19402\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__3738\ : LocalMux
    port map (
            O => \N__19399\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__3737\ : Odrv4
    port map (
            O => \N__19394\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__3736\ : LocalMux
    port map (
            O => \N__19391\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__3735\ : LocalMux
    port map (
            O => \N__19386\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__3734\ : InMux
    port map (
            O => \N__19369\,
            I => \N__19366\
        );

    \I__3733\ : LocalMux
    port map (
            O => \N__19366\,
            I => \N__19363\
        );

    \I__3732\ : Odrv4
    port map (
            O => \N__19363\,
            I => \uu2.bitmap_RNI1D952Z0Z_93\
        );

    \I__3731\ : InMux
    port map (
            O => \N__19360\,
            I => \N__19344\
        );

    \I__3730\ : InMux
    port map (
            O => \N__19359\,
            I => \N__19344\
        );

    \I__3729\ : InMux
    port map (
            O => \N__19358\,
            I => \N__19344\
        );

    \I__3728\ : InMux
    port map (
            O => \N__19357\,
            I => \N__19344\
        );

    \I__3727\ : InMux
    port map (
            O => \N__19356\,
            I => \N__19335\
        );

    \I__3726\ : InMux
    port map (
            O => \N__19355\,
            I => \N__19335\
        );

    \I__3725\ : InMux
    port map (
            O => \N__19354\,
            I => \N__19335\
        );

    \I__3724\ : InMux
    port map (
            O => \N__19353\,
            I => \N__19335\
        );

    \I__3723\ : LocalMux
    port map (
            O => \N__19344\,
            I => \Lab_UT.Sone_at_0\
        );

    \I__3722\ : LocalMux
    port map (
            O => \N__19335\,
            I => \Lab_UT.Sone_at_0\
        );

    \I__3721\ : CascadeMux
    port map (
            O => \N__19330\,
            I => \Lab_UT.Sone_at_0_cascade_\
        );

    \I__3720\ : InMux
    port map (
            O => \N__19327\,
            I => \N__19324\
        );

    \I__3719\ : LocalMux
    port map (
            O => \N__19324\,
            I => \N__19321\
        );

    \I__3718\ : Odrv4
    port map (
            O => \N__19321\,
            I => \Lab_UT.N_77_2\
        );

    \I__3717\ : CascadeMux
    port map (
            O => \N__19318\,
            I => \N__19312\
        );

    \I__3716\ : CascadeMux
    port map (
            O => \N__19317\,
            I => \N__19307\
        );

    \I__3715\ : CascadeMux
    port map (
            O => \N__19316\,
            I => \N__19301\
        );

    \I__3714\ : CascadeMux
    port map (
            O => \N__19315\,
            I => \N__19298\
        );

    \I__3713\ : InMux
    port map (
            O => \N__19312\,
            I => \N__19289\
        );

    \I__3712\ : InMux
    port map (
            O => \N__19311\,
            I => \N__19289\
        );

    \I__3711\ : InMux
    port map (
            O => \N__19310\,
            I => \N__19289\
        );

    \I__3710\ : InMux
    port map (
            O => \N__19307\,
            I => \N__19289\
        );

    \I__3709\ : InMux
    port map (
            O => \N__19306\,
            I => \N__19286\
        );

    \I__3708\ : InMux
    port map (
            O => \N__19305\,
            I => \N__19277\
        );

    \I__3707\ : InMux
    port map (
            O => \N__19304\,
            I => \N__19277\
        );

    \I__3706\ : InMux
    port map (
            O => \N__19301\,
            I => \N__19277\
        );

    \I__3705\ : InMux
    port map (
            O => \N__19298\,
            I => \N__19277\
        );

    \I__3704\ : LocalMux
    port map (
            O => \N__19289\,
            I => \Lab_UT.Sone_at_3\
        );

    \I__3703\ : LocalMux
    port map (
            O => \N__19286\,
            I => \Lab_UT.Sone_at_3\
        );

    \I__3702\ : LocalMux
    port map (
            O => \N__19277\,
            I => \Lab_UT.Sone_at_3\
        );

    \I__3701\ : InMux
    port map (
            O => \N__19270\,
            I => \N__19254\
        );

    \I__3700\ : InMux
    port map (
            O => \N__19269\,
            I => \N__19254\
        );

    \I__3699\ : InMux
    port map (
            O => \N__19268\,
            I => \N__19254\
        );

    \I__3698\ : InMux
    port map (
            O => \N__19267\,
            I => \N__19254\
        );

    \I__3697\ : InMux
    port map (
            O => \N__19266\,
            I => \N__19245\
        );

    \I__3696\ : InMux
    port map (
            O => \N__19265\,
            I => \N__19245\
        );

    \I__3695\ : InMux
    port map (
            O => \N__19264\,
            I => \N__19245\
        );

    \I__3694\ : InMux
    port map (
            O => \N__19263\,
            I => \N__19245\
        );

    \I__3693\ : LocalMux
    port map (
            O => \N__19254\,
            I => \Lab_UT.Sone_at_2\
        );

    \I__3692\ : LocalMux
    port map (
            O => \N__19245\,
            I => \Lab_UT.Sone_at_2\
        );

    \I__3691\ : InMux
    port map (
            O => \N__19240\,
            I => \N__19231\
        );

    \I__3690\ : InMux
    port map (
            O => \N__19239\,
            I => \N__19231\
        );

    \I__3689\ : InMux
    port map (
            O => \N__19238\,
            I => \N__19231\
        );

    \I__3688\ : LocalMux
    port map (
            O => \N__19231\,
            I => \resetGen.reset_countZ0Z_1\
        );

    \I__3687\ : InMux
    port map (
            O => \N__19228\,
            I => \N__19219\
        );

    \I__3686\ : InMux
    port map (
            O => \N__19227\,
            I => \N__19219\
        );

    \I__3685\ : InMux
    port map (
            O => \N__19226\,
            I => \N__19219\
        );

    \I__3684\ : LocalMux
    port map (
            O => \N__19219\,
            I => \N__19215\
        );

    \I__3683\ : InMux
    port map (
            O => \N__19218\,
            I => \N__19212\
        );

    \I__3682\ : Span4Mux_h
    port map (
            O => \N__19215\,
            I => \N__19209\
        );

    \I__3681\ : LocalMux
    port map (
            O => \N__19212\,
            I => \resetGen.reset_countZ0Z_0\
        );

    \I__3680\ : Odrv4
    port map (
            O => \N__19209\,
            I => \resetGen.reset_countZ0Z_0\
        );

    \I__3679\ : InMux
    port map (
            O => \N__19204\,
            I => \N__19201\
        );

    \I__3678\ : LocalMux
    port map (
            O => \N__19201\,
            I => \N__19198\
        );

    \I__3677\ : Span4Mux_h
    port map (
            O => \N__19198\,
            I => \N__19195\
        );

    \I__3676\ : Odrv4
    port map (
            O => \N__19195\,
            I => \resetGen.un241_ci\
        );

    \I__3675\ : CascadeMux
    port map (
            O => \N__19192\,
            I => \N__19188\
        );

    \I__3674\ : InMux
    port map (
            O => \N__19191\,
            I => \N__19183\
        );

    \I__3673\ : InMux
    port map (
            O => \N__19188\,
            I => \N__19176\
        );

    \I__3672\ : InMux
    port map (
            O => \N__19187\,
            I => \N__19176\
        );

    \I__3671\ : InMux
    port map (
            O => \N__19186\,
            I => \N__19176\
        );

    \I__3670\ : LocalMux
    port map (
            O => \N__19183\,
            I => \N__19173\
        );

    \I__3669\ : LocalMux
    port map (
            O => \N__19176\,
            I => \N__19168\
        );

    \I__3668\ : Span4Mux_v
    port map (
            O => \N__19173\,
            I => \N__19165\
        );

    \I__3667\ : InMux
    port map (
            O => \N__19172\,
            I => \N__19162\
        );

    \I__3666\ : InMux
    port map (
            O => \N__19171\,
            I => \N__19159\
        );

    \I__3665\ : Span4Mux_v
    port map (
            O => \N__19168\,
            I => \N__19154\
        );

    \I__3664\ : Span4Mux_v
    port map (
            O => \N__19165\,
            I => \N__19154\
        );

    \I__3663\ : LocalMux
    port map (
            O => \N__19162\,
            I => \resetGen.reset_countZ0Z_4\
        );

    \I__3662\ : LocalMux
    port map (
            O => \N__19159\,
            I => \resetGen.reset_countZ0Z_4\
        );

    \I__3661\ : Odrv4
    port map (
            O => \N__19154\,
            I => \resetGen.reset_countZ0Z_4\
        );

    \I__3660\ : CascadeMux
    port map (
            O => \N__19147\,
            I => \resetGen.un241_ci_cascade_\
        );

    \I__3659\ : InMux
    port map (
            O => \N__19144\,
            I => \N__19141\
        );

    \I__3658\ : LocalMux
    port map (
            O => \N__19141\,
            I => \N__19136\
        );

    \I__3657\ : InMux
    port map (
            O => \N__19140\,
            I => \N__19131\
        );

    \I__3656\ : InMux
    port map (
            O => \N__19139\,
            I => \N__19131\
        );

    \I__3655\ : Span4Mux_h
    port map (
            O => \N__19136\,
            I => \N__19128\
        );

    \I__3654\ : LocalMux
    port map (
            O => \N__19131\,
            I => \resetGen.reset_countZ0Z_2\
        );

    \I__3653\ : Odrv4
    port map (
            O => \N__19128\,
            I => \resetGen.reset_countZ0Z_2\
        );

    \I__3652\ : InMux
    port map (
            O => \N__19123\,
            I => \N__19120\
        );

    \I__3651\ : LocalMux
    port map (
            O => \N__19120\,
            I => \N__19117\
        );

    \I__3650\ : Span4Mux_v
    port map (
            O => \N__19117\,
            I => \N__19114\
        );

    \I__3649\ : Odrv4
    port map (
            O => \N__19114\,
            I => \Lab_UT.uu0.delay_lineZ0Z_1\
        );

    \I__3648\ : IoInMux
    port map (
            O => \N__19111\,
            I => \N__19108\
        );

    \I__3647\ : LocalMux
    port map (
            O => \N__19108\,
            I => \N__19105\
        );

    \I__3646\ : Span4Mux_s0_h
    port map (
            O => \N__19105\,
            I => \N__19102\
        );

    \I__3645\ : Span4Mux_h
    port map (
            O => \N__19102\,
            I => \N__19099\
        );

    \I__3644\ : Odrv4
    port map (
            O => \N__19099\,
            I => \Lab_UT.uu0.un11_l_count_i\
        );

    \I__3643\ : InMux
    port map (
            O => \N__19096\,
            I => \N__19093\
        );

    \I__3642\ : LocalMux
    port map (
            O => \N__19093\,
            I => \N__19090\
        );

    \I__3641\ : Odrv4
    port map (
            O => \N__19090\,
            I => \Lab_UT.L3_segment1_1_0_3\
        );

    \I__3640\ : CascadeMux
    port map (
            O => \N__19087\,
            I => \Lab_UT.L3_segment1_0_i_1_0_cascade_\
        );

    \I__3639\ : InMux
    port map (
            O => \N__19084\,
            I => \N__19081\
        );

    \I__3638\ : LocalMux
    port map (
            O => \N__19081\,
            I => \N__19078\
        );

    \I__3637\ : Odrv12
    port map (
            O => \N__19078\,
            I => \uu2.bitmapZ0Z_58\
        );

    \I__3636\ : InMux
    port map (
            O => \N__19075\,
            I => \N__19072\
        );

    \I__3635\ : LocalMux
    port map (
            O => \N__19072\,
            I => \Lab_UT.L3_segment1_0_i_1_1\
        );

    \I__3634\ : CascadeMux
    port map (
            O => \N__19069\,
            I => \N__19065\
        );

    \I__3633\ : InMux
    port map (
            O => \N__19068\,
            I => \N__19051\
        );

    \I__3632\ : InMux
    port map (
            O => \N__19065\,
            I => \N__19051\
        );

    \I__3631\ : InMux
    port map (
            O => \N__19064\,
            I => \N__19051\
        );

    \I__3630\ : InMux
    port map (
            O => \N__19063\,
            I => \N__19051\
        );

    \I__3629\ : InMux
    port map (
            O => \N__19062\,
            I => \N__19051\
        );

    \I__3628\ : LocalMux
    port map (
            O => \N__19051\,
            I => \N__19046\
        );

    \I__3627\ : InMux
    port map (
            O => \N__19050\,
            I => \N__19041\
        );

    \I__3626\ : InMux
    port map (
            O => \N__19049\,
            I => \N__19041\
        );

    \I__3625\ : Odrv4
    port map (
            O => \N__19046\,
            I => \uu2.w_addr_userZ0Z_0\
        );

    \I__3624\ : LocalMux
    port map (
            O => \N__19041\,
            I => \uu2.w_addr_userZ0Z_0\
        );

    \I__3623\ : CascadeMux
    port map (
            O => \N__19036\,
            I => \N__19031\
        );

    \I__3622\ : InMux
    port map (
            O => \N__19035\,
            I => \N__19027\
        );

    \I__3621\ : CascadeMux
    port map (
            O => \N__19034\,
            I => \N__19024\
        );

    \I__3620\ : InMux
    port map (
            O => \N__19031\,
            I => \N__19018\
        );

    \I__3619\ : InMux
    port map (
            O => \N__19030\,
            I => \N__19018\
        );

    \I__3618\ : LocalMux
    port map (
            O => \N__19027\,
            I => \N__19015\
        );

    \I__3617\ : InMux
    port map (
            O => \N__19024\,
            I => \N__19010\
        );

    \I__3616\ : InMux
    port map (
            O => \N__19023\,
            I => \N__19010\
        );

    \I__3615\ : LocalMux
    port map (
            O => \N__19018\,
            I => \N__19007\
        );

    \I__3614\ : Span4Mux_s3_v
    port map (
            O => \N__19015\,
            I => \N__19004\
        );

    \I__3613\ : LocalMux
    port map (
            O => \N__19010\,
            I => \uu2.w_addr_userZ0Z_2\
        );

    \I__3612\ : Odrv4
    port map (
            O => \N__19007\,
            I => \uu2.w_addr_userZ0Z_2\
        );

    \I__3611\ : Odrv4
    port map (
            O => \N__19004\,
            I => \uu2.w_addr_userZ0Z_2\
        );

    \I__3610\ : CascadeMux
    port map (
            O => \N__18997\,
            I => \N__18994\
        );

    \I__3609\ : InMux
    port map (
            O => \N__18994\,
            I => \N__18988\
        );

    \I__3608\ : InMux
    port map (
            O => \N__18993\,
            I => \N__18983\
        );

    \I__3607\ : InMux
    port map (
            O => \N__18992\,
            I => \N__18983\
        );

    \I__3606\ : InMux
    port map (
            O => \N__18991\,
            I => \N__18980\
        );

    \I__3605\ : LocalMux
    port map (
            O => \N__18988\,
            I => \uu2.w_addr_userZ0Z_3\
        );

    \I__3604\ : LocalMux
    port map (
            O => \N__18983\,
            I => \uu2.w_addr_userZ0Z_3\
        );

    \I__3603\ : LocalMux
    port map (
            O => \N__18980\,
            I => \uu2.w_addr_userZ0Z_3\
        );

    \I__3602\ : InMux
    port map (
            O => \N__18973\,
            I => \N__18970\
        );

    \I__3601\ : LocalMux
    port map (
            O => \N__18970\,
            I => \N__18964\
        );

    \I__3600\ : InMux
    port map (
            O => \N__18969\,
            I => \N__18955\
        );

    \I__3599\ : InMux
    port map (
            O => \N__18968\,
            I => \N__18955\
        );

    \I__3598\ : InMux
    port map (
            O => \N__18967\,
            I => \N__18955\
        );

    \I__3597\ : Span4Mux_h
    port map (
            O => \N__18964\,
            I => \N__18952\
        );

    \I__3596\ : InMux
    port map (
            O => \N__18963\,
            I => \N__18947\
        );

    \I__3595\ : InMux
    port map (
            O => \N__18962\,
            I => \N__18947\
        );

    \I__3594\ : LocalMux
    port map (
            O => \N__18955\,
            I => \uu2.w_addr_userZ0Z_1\
        );

    \I__3593\ : Odrv4
    port map (
            O => \N__18952\,
            I => \uu2.w_addr_userZ0Z_1\
        );

    \I__3592\ : LocalMux
    port map (
            O => \N__18947\,
            I => \uu2.w_addr_userZ0Z_1\
        );

    \I__3591\ : CascadeMux
    port map (
            O => \N__18940\,
            I => \resetGen.un252_ci_cascade_\
        );

    \I__3590\ : InMux
    port map (
            O => \N__18937\,
            I => \N__18934\
        );

    \I__3589\ : LocalMux
    port map (
            O => \N__18934\,
            I => \N__18930\
        );

    \I__3588\ : InMux
    port map (
            O => \N__18933\,
            I => \N__18927\
        );

    \I__3587\ : Span4Mux_v
    port map (
            O => \N__18930\,
            I => \N__18924\
        );

    \I__3586\ : LocalMux
    port map (
            O => \N__18927\,
            I => \resetGen.reset_countZ0Z_3\
        );

    \I__3585\ : Odrv4
    port map (
            O => \N__18924\,
            I => \resetGen.reset_countZ0Z_3\
        );

    \I__3584\ : CEMux
    port map (
            O => \N__18919\,
            I => \N__18915\
        );

    \I__3583\ : SRMux
    port map (
            O => \N__18918\,
            I => \N__18912\
        );

    \I__3582\ : LocalMux
    port map (
            O => \N__18915\,
            I => \N__18909\
        );

    \I__3581\ : LocalMux
    port map (
            O => \N__18912\,
            I => \N__18906\
        );

    \I__3580\ : Span4Mux_h
    port map (
            O => \N__18909\,
            I => \N__18903\
        );

    \I__3579\ : Odrv12
    port map (
            O => \N__18906\,
            I => \uu2.vram_wr_en_0_iZ0\
        );

    \I__3578\ : Odrv4
    port map (
            O => \N__18903\,
            I => \uu2.vram_wr_en_0_iZ0\
        );

    \I__3577\ : InMux
    port map (
            O => \N__18898\,
            I => \N__18895\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__18895\,
            I => \uu2.un1_w_user_lf_0\
        );

    \I__3575\ : CascadeMux
    port map (
            O => \N__18892\,
            I => \N__18888\
        );

    \I__3574\ : InMux
    port map (
            O => \N__18891\,
            I => \N__18883\
        );

    \I__3573\ : InMux
    port map (
            O => \N__18888\,
            I => \N__18883\
        );

    \I__3572\ : LocalMux
    port map (
            O => \N__18883\,
            I => \uu2.un3_w_addr_user\
        );

    \I__3571\ : InMux
    port map (
            O => \N__18880\,
            I => \N__18871\
        );

    \I__3570\ : InMux
    port map (
            O => \N__18879\,
            I => \N__18871\
        );

    \I__3569\ : InMux
    port map (
            O => \N__18878\,
            I => \N__18871\
        );

    \I__3568\ : LocalMux
    port map (
            O => \N__18871\,
            I => \uu2.un1_w_user_cr_0\
        );

    \I__3567\ : CascadeMux
    port map (
            O => \N__18868\,
            I => \uu2.un1_w_user_cr_0_cascade_\
        );

    \I__3566\ : InMux
    port map (
            O => \N__18865\,
            I => \N__18858\
        );

    \I__3565\ : InMux
    port map (
            O => \N__18864\,
            I => \N__18858\
        );

    \I__3564\ : InMux
    port map (
            O => \N__18863\,
            I => \N__18855\
        );

    \I__3563\ : LocalMux
    port map (
            O => \N__18858\,
            I => \N__18852\
        );

    \I__3562\ : LocalMux
    port map (
            O => \N__18855\,
            I => \uu2.N_71\
        );

    \I__3561\ : Odrv12
    port map (
            O => \N__18852\,
            I => \uu2.N_71\
        );

    \I__3560\ : CascadeMux
    port map (
            O => \N__18847\,
            I => \uu2.un4_w_user_data_rdyZ0Z_0_cascade_\
        );

    \I__3559\ : InMux
    port map (
            O => \N__18844\,
            I => \N__18841\
        );

    \I__3558\ : LocalMux
    port map (
            O => \N__18841\,
            I => \N__18838\
        );

    \I__3557\ : Span4Mux_s3_h
    port map (
            O => \N__18838\,
            I => \N__18835\
        );

    \I__3556\ : Span4Mux_h
    port map (
            O => \N__18835\,
            I => \N__18832\
        );

    \I__3555\ : Odrv4
    port map (
            O => \N__18832\,
            I => \uu2.mem0.w_data_6\
        );

    \I__3554\ : InMux
    port map (
            O => \N__18829\,
            I => \N__18826\
        );

    \I__3553\ : LocalMux
    port map (
            O => \N__18826\,
            I => \uu2.un1_w_user_crZ0Z_4\
        );

    \I__3552\ : InMux
    port map (
            O => \N__18823\,
            I => \N__18820\
        );

    \I__3551\ : LocalMux
    port map (
            O => \N__18820\,
            I => \uu2.un1_w_user_lfZ0Z_4\
        );

    \I__3550\ : InMux
    port map (
            O => \N__18817\,
            I => \N__18814\
        );

    \I__3549\ : LocalMux
    port map (
            O => \N__18814\,
            I => \N__18811\
        );

    \I__3548\ : Span4Mux_s3_h
    port map (
            O => \N__18811\,
            I => \N__18808\
        );

    \I__3547\ : Span4Mux_h
    port map (
            O => \N__18808\,
            I => \N__18805\
        );

    \I__3546\ : Odrv4
    port map (
            O => \N__18805\,
            I => \uu2.mem0.w_data_2\
        );

    \I__3545\ : InMux
    port map (
            O => \N__18802\,
            I => \N__18787\
        );

    \I__3544\ : InMux
    port map (
            O => \N__18801\,
            I => \N__18787\
        );

    \I__3543\ : InMux
    port map (
            O => \N__18800\,
            I => \N__18787\
        );

    \I__3542\ : InMux
    port map (
            O => \N__18799\,
            I => \N__18787\
        );

    \I__3541\ : InMux
    port map (
            O => \N__18798\,
            I => \N__18787\
        );

    \I__3540\ : LocalMux
    port map (
            O => \N__18787\,
            I => \N__18782\
        );

    \I__3539\ : InMux
    port map (
            O => \N__18786\,
            I => \N__18779\
        );

    \I__3538\ : InMux
    port map (
            O => \N__18785\,
            I => \N__18776\
        );

    \I__3537\ : Span4Mux_v
    port map (
            O => \N__18782\,
            I => \N__18764\
        );

    \I__3536\ : LocalMux
    port map (
            O => \N__18779\,
            I => \N__18764\
        );

    \I__3535\ : LocalMux
    port map (
            O => \N__18776\,
            I => \N__18764\
        );

    \I__3534\ : InMux
    port map (
            O => \N__18775\,
            I => \N__18761\
        );

    \I__3533\ : InMux
    port map (
            O => \N__18774\,
            I => \N__18752\
        );

    \I__3532\ : InMux
    port map (
            O => \N__18773\,
            I => \N__18752\
        );

    \I__3531\ : InMux
    port map (
            O => \N__18772\,
            I => \N__18752\
        );

    \I__3530\ : InMux
    port map (
            O => \N__18771\,
            I => \N__18752\
        );

    \I__3529\ : Span4Mux_h
    port map (
            O => \N__18764\,
            I => \N__18745\
        );

    \I__3528\ : LocalMux
    port map (
            O => \N__18761\,
            I => \N__18742\
        );

    \I__3527\ : LocalMux
    port map (
            O => \N__18752\,
            I => \N__18739\
        );

    \I__3526\ : InMux
    port map (
            O => \N__18751\,
            I => \N__18734\
        );

    \I__3525\ : InMux
    port map (
            O => \N__18750\,
            I => \N__18734\
        );

    \I__3524\ : InMux
    port map (
            O => \N__18749\,
            I => \N__18731\
        );

    \I__3523\ : InMux
    port map (
            O => \N__18748\,
            I => \N__18728\
        );

    \I__3522\ : Odrv4
    port map (
            O => \N__18745\,
            I => \uu2.un4_w_user_data_rdyZ0Z_0\
        );

    \I__3521\ : Odrv12
    port map (
            O => \N__18742\,
            I => \uu2.un4_w_user_data_rdyZ0Z_0\
        );

    \I__3520\ : Odrv4
    port map (
            O => \N__18739\,
            I => \uu2.un4_w_user_data_rdyZ0Z_0\
        );

    \I__3519\ : LocalMux
    port map (
            O => \N__18734\,
            I => \uu2.un4_w_user_data_rdyZ0Z_0\
        );

    \I__3518\ : LocalMux
    port map (
            O => \N__18731\,
            I => \uu2.un4_w_user_data_rdyZ0Z_0\
        );

    \I__3517\ : LocalMux
    port map (
            O => \N__18728\,
            I => \uu2.un4_w_user_data_rdyZ0Z_0\
        );

    \I__3516\ : CascadeMux
    port map (
            O => \N__18715\,
            I => \N__18712\
        );

    \I__3515\ : InMux
    port map (
            O => \N__18712\,
            I => \N__18709\
        );

    \I__3514\ : LocalMux
    port map (
            O => \N__18709\,
            I => \N__18706\
        );

    \I__3513\ : Span12Mux_s7_h
    port map (
            O => \N__18706\,
            I => \N__18703\
        );

    \I__3512\ : Odrv12
    port map (
            O => \N__18703\,
            I => \uu2.mem0.w_addr_0\
        );

    \I__3511\ : CascadeMux
    port map (
            O => \N__18700\,
            I => \Lab_UT.uu0.un4_l_count_14_cascade_\
        );

    \I__3510\ : CascadeMux
    port map (
            O => \N__18697\,
            I => \Lab_UT.uu0.un187_ci_1_cascade_\
        );

    \I__3509\ : CascadeMux
    port map (
            O => \N__18694\,
            I => \N__18691\
        );

    \I__3508\ : InMux
    port map (
            O => \N__18691\,
            I => \N__18685\
        );

    \I__3507\ : InMux
    port map (
            O => \N__18690\,
            I => \N__18678\
        );

    \I__3506\ : InMux
    port map (
            O => \N__18689\,
            I => \N__18678\
        );

    \I__3505\ : InMux
    port map (
            O => \N__18688\,
            I => \N__18678\
        );

    \I__3504\ : LocalMux
    port map (
            O => \N__18685\,
            I => \Lab_UT.uu0.un154_ci_9\
        );

    \I__3503\ : LocalMux
    port map (
            O => \N__18678\,
            I => \Lab_UT.uu0.un154_ci_9\
        );

    \I__3502\ : CascadeMux
    port map (
            O => \N__18673\,
            I => \N__18667\
        );

    \I__3501\ : CascadeMux
    port map (
            O => \N__18672\,
            I => \N__18664\
        );

    \I__3500\ : CascadeMux
    port map (
            O => \N__18671\,
            I => \N__18661\
        );

    \I__3499\ : InMux
    port map (
            O => \N__18670\,
            I => \N__18656\
        );

    \I__3498\ : InMux
    port map (
            O => \N__18667\,
            I => \N__18656\
        );

    \I__3497\ : InMux
    port map (
            O => \N__18664\,
            I => \N__18651\
        );

    \I__3496\ : InMux
    port map (
            O => \N__18661\,
            I => \N__18651\
        );

    \I__3495\ : LocalMux
    port map (
            O => \N__18656\,
            I => \Lab_UT.uu0.l_countZ0Z_14\
        );

    \I__3494\ : LocalMux
    port map (
            O => \N__18651\,
            I => \Lab_UT.uu0.l_countZ0Z_14\
        );

    \I__3493\ : InMux
    port map (
            O => \N__18646\,
            I => \N__18640\
        );

    \I__3492\ : InMux
    port map (
            O => \N__18645\,
            I => \N__18633\
        );

    \I__3491\ : InMux
    port map (
            O => \N__18644\,
            I => \N__18633\
        );

    \I__3490\ : InMux
    port map (
            O => \N__18643\,
            I => \N__18633\
        );

    \I__3489\ : LocalMux
    port map (
            O => \N__18640\,
            I => \N__18628\
        );

    \I__3488\ : LocalMux
    port map (
            O => \N__18633\,
            I => \N__18628\
        );

    \I__3487\ : Span4Mux_h
    port map (
            O => \N__18628\,
            I => \N__18625\
        );

    \I__3486\ : Odrv4
    port map (
            O => \N__18625\,
            I => \Lab_UT.uu0.un4_l_count_0_8\
        );

    \I__3485\ : InMux
    port map (
            O => \N__18622\,
            I => \N__18613\
        );

    \I__3484\ : InMux
    port map (
            O => \N__18621\,
            I => \N__18613\
        );

    \I__3483\ : InMux
    port map (
            O => \N__18620\,
            I => \N__18613\
        );

    \I__3482\ : LocalMux
    port map (
            O => \N__18613\,
            I => \Lab_UT.uu0.un198_ci_2\
        );

    \I__3481\ : CascadeMux
    port map (
            O => \N__18610\,
            I => \N__18605\
        );

    \I__3480\ : CascadeMux
    port map (
            O => \N__18609\,
            I => \N__18598\
        );

    \I__3479\ : CascadeMux
    port map (
            O => \N__18608\,
            I => \N__18595\
        );

    \I__3478\ : InMux
    port map (
            O => \N__18605\,
            I => \N__18585\
        );

    \I__3477\ : InMux
    port map (
            O => \N__18604\,
            I => \N__18585\
        );

    \I__3476\ : InMux
    port map (
            O => \N__18603\,
            I => \N__18585\
        );

    \I__3475\ : InMux
    port map (
            O => \N__18602\,
            I => \N__18582\
        );

    \I__3474\ : InMux
    port map (
            O => \N__18601\,
            I => \N__18577\
        );

    \I__3473\ : InMux
    port map (
            O => \N__18598\,
            I => \N__18577\
        );

    \I__3472\ : InMux
    port map (
            O => \N__18595\,
            I => \N__18568\
        );

    \I__3471\ : InMux
    port map (
            O => \N__18594\,
            I => \N__18568\
        );

    \I__3470\ : InMux
    port map (
            O => \N__18593\,
            I => \N__18568\
        );

    \I__3469\ : InMux
    port map (
            O => \N__18592\,
            I => \N__18568\
        );

    \I__3468\ : LocalMux
    port map (
            O => \N__18585\,
            I => \Lab_UT.uu0.un110_ci\
        );

    \I__3467\ : LocalMux
    port map (
            O => \N__18582\,
            I => \Lab_UT.uu0.un110_ci\
        );

    \I__3466\ : LocalMux
    port map (
            O => \N__18577\,
            I => \Lab_UT.uu0.un110_ci\
        );

    \I__3465\ : LocalMux
    port map (
            O => \N__18568\,
            I => \Lab_UT.uu0.un110_ci\
        );

    \I__3464\ : InMux
    port map (
            O => \N__18559\,
            I => \N__18547\
        );

    \I__3463\ : InMux
    port map (
            O => \N__18558\,
            I => \N__18547\
        );

    \I__3462\ : InMux
    port map (
            O => \N__18557\,
            I => \N__18547\
        );

    \I__3461\ : InMux
    port map (
            O => \N__18556\,
            I => \N__18540\
        );

    \I__3460\ : InMux
    port map (
            O => \N__18555\,
            I => \N__18540\
        );

    \I__3459\ : InMux
    port map (
            O => \N__18554\,
            I => \N__18540\
        );

    \I__3458\ : LocalMux
    port map (
            O => \N__18547\,
            I => \Lab_UT.uu0.l_countZ0Z_8\
        );

    \I__3457\ : LocalMux
    port map (
            O => \N__18540\,
            I => \Lab_UT.uu0.l_countZ0Z_8\
        );

    \I__3456\ : CEMux
    port map (
            O => \N__18535\,
            I => \N__18532\
        );

    \I__3455\ : LocalMux
    port map (
            O => \N__18532\,
            I => \N__18529\
        );

    \I__3454\ : Span4Mux_s2_v
    port map (
            O => \N__18529\,
            I => \N__18526\
        );

    \I__3453\ : Odrv4
    port map (
            O => \N__18526\,
            I => \uu2.un28_w_addr_user_i_0\
        );

    \I__3452\ : CascadeMux
    port map (
            O => \N__18523\,
            I => \uu2.un1_w_user_lf_0_cascade_\
        );

    \I__3451\ : CascadeMux
    port map (
            O => \N__18520\,
            I => \Lab_UT.uu0.un99_ci_0_cascade_\
        );

    \I__3450\ : CascadeMux
    port map (
            O => \N__18517\,
            I => \N__18514\
        );

    \I__3449\ : InMux
    port map (
            O => \N__18514\,
            I => \N__18508\
        );

    \I__3448\ : InMux
    port map (
            O => \N__18513\,
            I => \N__18508\
        );

    \I__3447\ : LocalMux
    port map (
            O => \N__18508\,
            I => \Lab_UT.uu0.un88_ci_3\
        );

    \I__3446\ : CascadeMux
    port map (
            O => \N__18505\,
            I => \Lab_UT.uu0.un88_ci_3_cascade_\
        );

    \I__3445\ : InMux
    port map (
            O => \N__18502\,
            I => \N__18495\
        );

    \I__3444\ : InMux
    port map (
            O => \N__18501\,
            I => \N__18495\
        );

    \I__3443\ : InMux
    port map (
            O => \N__18500\,
            I => \N__18492\
        );

    \I__3442\ : LocalMux
    port map (
            O => \N__18495\,
            I => \Lab_UT.uu0.l_countZ0Z_7\
        );

    \I__3441\ : LocalMux
    port map (
            O => \N__18492\,
            I => \Lab_UT.uu0.l_countZ0Z_7\
        );

    \I__3440\ : CascadeMux
    port map (
            O => \N__18487\,
            I => \N__18483\
        );

    \I__3439\ : CascadeMux
    port map (
            O => \N__18486\,
            I => \N__18480\
        );

    \I__3438\ : InMux
    port map (
            O => \N__18483\,
            I => \N__18476\
        );

    \I__3437\ : InMux
    port map (
            O => \N__18480\,
            I => \N__18471\
        );

    \I__3436\ : InMux
    port map (
            O => \N__18479\,
            I => \N__18471\
        );

    \I__3435\ : LocalMux
    port map (
            O => \N__18476\,
            I => \N__18468\
        );

    \I__3434\ : LocalMux
    port map (
            O => \N__18471\,
            I => \Lab_UT.uu0.l_countZ0Z_17\
        );

    \I__3433\ : Odrv4
    port map (
            O => \N__18468\,
            I => \Lab_UT.uu0.l_countZ0Z_17\
        );

    \I__3432\ : CascadeMux
    port map (
            O => \N__18463\,
            I => \Lab_UT.uu0.un110_ci_cascade_\
        );

    \I__3431\ : InMux
    port map (
            O => \N__18460\,
            I => \N__18457\
        );

    \I__3430\ : LocalMux
    port map (
            O => \N__18457\,
            I => \Lab_UT.uu0.un220_ci\
        );

    \I__3429\ : InMux
    port map (
            O => \N__18454\,
            I => \N__18447\
        );

    \I__3428\ : InMux
    port map (
            O => \N__18453\,
            I => \N__18440\
        );

    \I__3427\ : InMux
    port map (
            O => \N__18452\,
            I => \N__18440\
        );

    \I__3426\ : InMux
    port map (
            O => \N__18451\,
            I => \N__18440\
        );

    \I__3425\ : InMux
    port map (
            O => \N__18450\,
            I => \N__18437\
        );

    \I__3424\ : LocalMux
    port map (
            O => \N__18447\,
            I => \Lab_UT.uu0.l_countZ0Z_9\
        );

    \I__3423\ : LocalMux
    port map (
            O => \N__18440\,
            I => \Lab_UT.uu0.l_countZ0Z_9\
        );

    \I__3422\ : LocalMux
    port map (
            O => \N__18437\,
            I => \Lab_UT.uu0.l_countZ0Z_9\
        );

    \I__3421\ : InMux
    port map (
            O => \N__18430\,
            I => \N__18424\
        );

    \I__3420\ : InMux
    port map (
            O => \N__18429\,
            I => \N__18421\
        );

    \I__3419\ : InMux
    port map (
            O => \N__18428\,
            I => \N__18416\
        );

    \I__3418\ : InMux
    port map (
            O => \N__18427\,
            I => \N__18416\
        );

    \I__3417\ : LocalMux
    port map (
            O => \N__18424\,
            I => \Lab_UT.uu0.l_countZ0Z_10\
        );

    \I__3416\ : LocalMux
    port map (
            O => \N__18421\,
            I => \Lab_UT.uu0.l_countZ0Z_10\
        );

    \I__3415\ : LocalMux
    port map (
            O => \N__18416\,
            I => \Lab_UT.uu0.l_countZ0Z_10\
        );

    \I__3414\ : InMux
    port map (
            O => \N__18409\,
            I => \N__18406\
        );

    \I__3413\ : LocalMux
    port map (
            O => \N__18406\,
            I => \N__18403\
        );

    \I__3412\ : Odrv4
    port map (
            O => \N__18403\,
            I => \Lab_UT.dictrl.decoder.g0_3Z0Z_0\
        );

    \I__3411\ : CascadeMux
    port map (
            O => \N__18400\,
            I => \N__18397\
        );

    \I__3410\ : InMux
    port map (
            O => \N__18397\,
            I => \N__18394\
        );

    \I__3409\ : LocalMux
    port map (
            O => \N__18394\,
            I => \N__18391\
        );

    \I__3408\ : Span4Mux_h
    port map (
            O => \N__18391\,
            I => \N__18388\
        );

    \I__3407\ : Odrv4
    port map (
            O => \N__18388\,
            I => \Lab_UT.dictrl.de_cr_1_2\
        );

    \I__3406\ : InMux
    port map (
            O => \N__18385\,
            I => \N__18382\
        );

    \I__3405\ : LocalMux
    port map (
            O => \N__18382\,
            I => \Lab_UT.dictrl.decoder.g0_4Z0Z_3\
        );

    \I__3404\ : CascadeMux
    port map (
            O => \N__18379\,
            I => \Lab_UT.dictrl.decoder.g0_3_2_cascade_\
        );

    \I__3403\ : CascadeMux
    port map (
            O => \N__18376\,
            I => \N__18372\
        );

    \I__3402\ : InMux
    port map (
            O => \N__18375\,
            I => \N__18368\
        );

    \I__3401\ : InMux
    port map (
            O => \N__18372\,
            I => \N__18361\
        );

    \I__3400\ : InMux
    port map (
            O => \N__18371\,
            I => \N__18361\
        );

    \I__3399\ : LocalMux
    port map (
            O => \N__18368\,
            I => \N__18358\
        );

    \I__3398\ : InMux
    port map (
            O => \N__18367\,
            I => \N__18353\
        );

    \I__3397\ : InMux
    port map (
            O => \N__18366\,
            I => \N__18353\
        );

    \I__3396\ : LocalMux
    port map (
            O => \N__18361\,
            I => \N__18348\
        );

    \I__3395\ : Span4Mux_h
    port map (
            O => \N__18358\,
            I => \N__18348\
        );

    \I__3394\ : LocalMux
    port map (
            O => \N__18353\,
            I => \Lab_UT_dictrl_decoder_de_cr_1_1\
        );

    \I__3393\ : Odrv4
    port map (
            O => \N__18348\,
            I => \Lab_UT_dictrl_decoder_de_cr_1_1\
        );

    \I__3392\ : CascadeMux
    port map (
            O => \N__18343\,
            I => \N__18340\
        );

    \I__3391\ : InMux
    port map (
            O => \N__18340\,
            I => \N__18337\
        );

    \I__3390\ : LocalMux
    port map (
            O => \N__18337\,
            I => \N__18334\
        );

    \I__3389\ : Odrv4
    port map (
            O => \N__18334\,
            I => \Lab_UT.dictrl.de_cr_2_0\
        );

    \I__3388\ : CascadeMux
    port map (
            O => \N__18331\,
            I => \N__18328\
        );

    \I__3387\ : InMux
    port map (
            O => \N__18328\,
            I => \N__18325\
        );

    \I__3386\ : LocalMux
    port map (
            O => \N__18325\,
            I => \Lab_UT.dictrl.decoder.g0_4_1\
        );

    \I__3385\ : CascadeMux
    port map (
            O => \N__18322\,
            I => \N__18314\
        );

    \I__3384\ : CascadeMux
    port map (
            O => \N__18321\,
            I => \N__18311\
        );

    \I__3383\ : CascadeMux
    port map (
            O => \N__18320\,
            I => \N__18308\
        );

    \I__3382\ : InMux
    port map (
            O => \N__18319\,
            I => \N__18301\
        );

    \I__3381\ : InMux
    port map (
            O => \N__18318\,
            I => \N__18301\
        );

    \I__3380\ : InMux
    port map (
            O => \N__18317\,
            I => \N__18294\
        );

    \I__3379\ : InMux
    port map (
            O => \N__18314\,
            I => \N__18294\
        );

    \I__3378\ : InMux
    port map (
            O => \N__18311\,
            I => \N__18294\
        );

    \I__3377\ : InMux
    port map (
            O => \N__18308\,
            I => \N__18287\
        );

    \I__3376\ : InMux
    port map (
            O => \N__18307\,
            I => \N__18287\
        );

    \I__3375\ : InMux
    port map (
            O => \N__18306\,
            I => \N__18287\
        );

    \I__3374\ : LocalMux
    port map (
            O => \N__18301\,
            I => \buart__rx_bitcount_4\
        );

    \I__3373\ : LocalMux
    port map (
            O => \N__18294\,
            I => \buart__rx_bitcount_4\
        );

    \I__3372\ : LocalMux
    port map (
            O => \N__18287\,
            I => \buart__rx_bitcount_4\
        );

    \I__3371\ : InMux
    port map (
            O => \N__18280\,
            I => \N__18275\
        );

    \I__3370\ : InMux
    port map (
            O => \N__18279\,
            I => \N__18264\
        );

    \I__3369\ : InMux
    port map (
            O => \N__18278\,
            I => \N__18264\
        );

    \I__3368\ : LocalMux
    port map (
            O => \N__18275\,
            I => \N__18261\
        );

    \I__3367\ : InMux
    port map (
            O => \N__18274\,
            I => \N__18254\
        );

    \I__3366\ : InMux
    port map (
            O => \N__18273\,
            I => \N__18254\
        );

    \I__3365\ : InMux
    port map (
            O => \N__18272\,
            I => \N__18254\
        );

    \I__3364\ : InMux
    port map (
            O => \N__18271\,
            I => \N__18247\
        );

    \I__3363\ : InMux
    port map (
            O => \N__18270\,
            I => \N__18247\
        );

    \I__3362\ : InMux
    port map (
            O => \N__18269\,
            I => \N__18247\
        );

    \I__3361\ : LocalMux
    port map (
            O => \N__18264\,
            I => \buart__rx_bitcount_3\
        );

    \I__3360\ : Odrv4
    port map (
            O => \N__18261\,
            I => \buart__rx_bitcount_3\
        );

    \I__3359\ : LocalMux
    port map (
            O => \N__18254\,
            I => \buart__rx_bitcount_3\
        );

    \I__3358\ : LocalMux
    port map (
            O => \N__18247\,
            I => \buart__rx_bitcount_3\
        );

    \I__3357\ : InMux
    port map (
            O => \N__18238\,
            I => \N__18227\
        );

    \I__3356\ : InMux
    port map (
            O => \N__18237\,
            I => \N__18227\
        );

    \I__3355\ : InMux
    port map (
            O => \N__18236\,
            I => \N__18217\
        );

    \I__3354\ : InMux
    port map (
            O => \N__18235\,
            I => \N__18217\
        );

    \I__3353\ : InMux
    port map (
            O => \N__18234\,
            I => \N__18217\
        );

    \I__3352\ : InMux
    port map (
            O => \N__18233\,
            I => \N__18212\
        );

    \I__3351\ : InMux
    port map (
            O => \N__18232\,
            I => \N__18212\
        );

    \I__3350\ : LocalMux
    port map (
            O => \N__18227\,
            I => \N__18209\
        );

    \I__3349\ : InMux
    port map (
            O => \N__18226\,
            I => \N__18204\
        );

    \I__3348\ : InMux
    port map (
            O => \N__18225\,
            I => \N__18204\
        );

    \I__3347\ : InMux
    port map (
            O => \N__18224\,
            I => \N__18201\
        );

    \I__3346\ : LocalMux
    port map (
            O => \N__18217\,
            I => \buart__rx_bitcount_2\
        );

    \I__3345\ : LocalMux
    port map (
            O => \N__18212\,
            I => \buart__rx_bitcount_2\
        );

    \I__3344\ : Odrv4
    port map (
            O => \N__18209\,
            I => \buart__rx_bitcount_2\
        );

    \I__3343\ : LocalMux
    port map (
            O => \N__18204\,
            I => \buart__rx_bitcount_2\
        );

    \I__3342\ : LocalMux
    port map (
            O => \N__18201\,
            I => \buart__rx_bitcount_2\
        );

    \I__3341\ : CascadeMux
    port map (
            O => \N__18190\,
            I => \Lab_UT.dictrl.g0_8_cascade_\
        );

    \I__3340\ : InMux
    port map (
            O => \N__18187\,
            I => \N__18183\
        );

    \I__3339\ : CascadeMux
    port map (
            O => \N__18186\,
            I => \N__18180\
        );

    \I__3338\ : LocalMux
    port map (
            O => \N__18183\,
            I => \N__18176\
        );

    \I__3337\ : InMux
    port map (
            O => \N__18180\,
            I => \N__18168\
        );

    \I__3336\ : InMux
    port map (
            O => \N__18179\,
            I => \N__18165\
        );

    \I__3335\ : Span4Mux_v
    port map (
            O => \N__18176\,
            I => \N__18162\
        );

    \I__3334\ : InMux
    port map (
            O => \N__18175\,
            I => \N__18155\
        );

    \I__3333\ : InMux
    port map (
            O => \N__18174\,
            I => \N__18155\
        );

    \I__3332\ : InMux
    port map (
            O => \N__18173\,
            I => \N__18155\
        );

    \I__3331\ : InMux
    port map (
            O => \N__18172\,
            I => \N__18152\
        );

    \I__3330\ : InMux
    port map (
            O => \N__18171\,
            I => \N__18149\
        );

    \I__3329\ : LocalMux
    port map (
            O => \N__18168\,
            I => \N__18146\
        );

    \I__3328\ : LocalMux
    port map (
            O => \N__18165\,
            I => \N__18143\
        );

    \I__3327\ : Odrv4
    port map (
            O => \N__18162\,
            I => \buart__rx_valid_2_0\
        );

    \I__3326\ : LocalMux
    port map (
            O => \N__18155\,
            I => \buart__rx_valid_2_0\
        );

    \I__3325\ : LocalMux
    port map (
            O => \N__18152\,
            I => \buart__rx_valid_2_0\
        );

    \I__3324\ : LocalMux
    port map (
            O => \N__18149\,
            I => \buart__rx_valid_2_0\
        );

    \I__3323\ : Odrv4
    port map (
            O => \N__18146\,
            I => \buart__rx_valid_2_0\
        );

    \I__3322\ : Odrv4
    port map (
            O => \N__18143\,
            I => \buart__rx_valid_2_0\
        );

    \I__3321\ : InMux
    port map (
            O => \N__18130\,
            I => \N__18127\
        );

    \I__3320\ : LocalMux
    port map (
            O => \N__18127\,
            I => \N__18124\
        );

    \I__3319\ : Span4Mux_h
    port map (
            O => \N__18124\,
            I => \N__18121\
        );

    \I__3318\ : Span4Mux_v
    port map (
            O => \N__18121\,
            I => \N__18118\
        );

    \I__3317\ : Odrv4
    port map (
            O => \N__18118\,
            I => \Lab_UT.dictrl.g0_11\
        );

    \I__3316\ : InMux
    port map (
            O => \N__18115\,
            I => \N__18112\
        );

    \I__3315\ : LocalMux
    port map (
            O => \N__18112\,
            I => \N__18108\
        );

    \I__3314\ : InMux
    port map (
            O => \N__18111\,
            I => \N__18105\
        );

    \I__3313\ : Span4Mux_v
    port map (
            O => \N__18108\,
            I => \N__18102\
        );

    \I__3312\ : LocalMux
    port map (
            O => \N__18105\,
            I => \N__18099\
        );

    \I__3311\ : Span4Mux_h
    port map (
            O => \N__18102\,
            I => \N__18096\
        );

    \I__3310\ : Span4Mux_h
    port map (
            O => \N__18099\,
            I => \N__18093\
        );

    \I__3309\ : Odrv4
    port map (
            O => \N__18096\,
            I => \Lab_UT.dictrl.currState_2_RNIEPCJZ0Z_1\
        );

    \I__3308\ : Odrv4
    port map (
            O => \N__18093\,
            I => \Lab_UT.dictrl.currState_2_RNIEPCJZ0Z_1\
        );

    \I__3307\ : InMux
    port map (
            O => \N__18088\,
            I => \N__18085\
        );

    \I__3306\ : LocalMux
    port map (
            O => \N__18085\,
            I => \N__18081\
        );

    \I__3305\ : InMux
    port map (
            O => \N__18084\,
            I => \N__18078\
        );

    \I__3304\ : Span4Mux_h
    port map (
            O => \N__18081\,
            I => \N__18075\
        );

    \I__3303\ : LocalMux
    port map (
            O => \N__18078\,
            I => \Lab_UT.dictrl.nextState_0_3\
        );

    \I__3302\ : Odrv4
    port map (
            O => \N__18075\,
            I => \Lab_UT.dictrl.nextState_0_3\
        );

    \I__3301\ : InMux
    port map (
            O => \N__18070\,
            I => \N__18067\
        );

    \I__3300\ : LocalMux
    port map (
            O => \N__18067\,
            I => \Lab_UT.dictrl.N_1612_0\
        );

    \I__3299\ : InMux
    port map (
            O => \N__18064\,
            I => \N__18048\
        );

    \I__3298\ : InMux
    port map (
            O => \N__18063\,
            I => \N__18048\
        );

    \I__3297\ : InMux
    port map (
            O => \N__18062\,
            I => \N__18043\
        );

    \I__3296\ : InMux
    port map (
            O => \N__18061\,
            I => \N__18038\
        );

    \I__3295\ : InMux
    port map (
            O => \N__18060\,
            I => \N__18031\
        );

    \I__3294\ : InMux
    port map (
            O => \N__18059\,
            I => \N__18031\
        );

    \I__3293\ : InMux
    port map (
            O => \N__18058\,
            I => \N__18031\
        );

    \I__3292\ : InMux
    port map (
            O => \N__18057\,
            I => \N__18026\
        );

    \I__3291\ : InMux
    port map (
            O => \N__18056\,
            I => \N__18026\
        );

    \I__3290\ : InMux
    port map (
            O => \N__18055\,
            I => \N__18023\
        );

    \I__3289\ : InMux
    port map (
            O => \N__18054\,
            I => \N__18018\
        );

    \I__3288\ : InMux
    port map (
            O => \N__18053\,
            I => \N__18018\
        );

    \I__3287\ : LocalMux
    port map (
            O => \N__18048\,
            I => \N__18015\
        );

    \I__3286\ : CascadeMux
    port map (
            O => \N__18047\,
            I => \N__18010\
        );

    \I__3285\ : InMux
    port map (
            O => \N__18046\,
            I => \N__18003\
        );

    \I__3284\ : LocalMux
    port map (
            O => \N__18043\,
            I => \N__18000\
        );

    \I__3283\ : InMux
    port map (
            O => \N__18042\,
            I => \N__17997\
        );

    \I__3282\ : InMux
    port map (
            O => \N__18041\,
            I => \N__17994\
        );

    \I__3281\ : LocalMux
    port map (
            O => \N__18038\,
            I => \N__17987\
        );

    \I__3280\ : LocalMux
    port map (
            O => \N__18031\,
            I => \N__17987\
        );

    \I__3279\ : LocalMux
    port map (
            O => \N__18026\,
            I => \N__17987\
        );

    \I__3278\ : LocalMux
    port map (
            O => \N__18023\,
            I => \N__17982\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__18018\,
            I => \N__17982\
        );

    \I__3276\ : Span4Mux_v
    port map (
            O => \N__18015\,
            I => \N__17979\
        );

    \I__3275\ : InMux
    port map (
            O => \N__18014\,
            I => \N__17976\
        );

    \I__3274\ : InMux
    port map (
            O => \N__18013\,
            I => \N__17973\
        );

    \I__3273\ : InMux
    port map (
            O => \N__18010\,
            I => \N__17966\
        );

    \I__3272\ : InMux
    port map (
            O => \N__18009\,
            I => \N__17966\
        );

    \I__3271\ : InMux
    port map (
            O => \N__18008\,
            I => \N__17966\
        );

    \I__3270\ : InMux
    port map (
            O => \N__18007\,
            I => \N__17963\
        );

    \I__3269\ : InMux
    port map (
            O => \N__18006\,
            I => \N__17960\
        );

    \I__3268\ : LocalMux
    port map (
            O => \N__18003\,
            I => \N__17951\
        );

    \I__3267\ : Span4Mux_h
    port map (
            O => \N__18000\,
            I => \N__17951\
        );

    \I__3266\ : LocalMux
    port map (
            O => \N__17997\,
            I => \N__17951\
        );

    \I__3265\ : LocalMux
    port map (
            O => \N__17994\,
            I => \N__17951\
        );

    \I__3264\ : Span4Mux_v
    port map (
            O => \N__17987\,
            I => \N__17946\
        );

    \I__3263\ : Span4Mux_v
    port map (
            O => \N__17982\,
            I => \N__17946\
        );

    \I__3262\ : Odrv4
    port map (
            O => \N__17979\,
            I => \Lab_UT.dictrl.currState_2_RNI2P2AZ0Z_2\
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__17976\,
            I => \Lab_UT.dictrl.currState_2_RNI2P2AZ0Z_2\
        );

    \I__3260\ : LocalMux
    port map (
            O => \N__17973\,
            I => \Lab_UT.dictrl.currState_2_RNI2P2AZ0Z_2\
        );

    \I__3259\ : LocalMux
    port map (
            O => \N__17966\,
            I => \Lab_UT.dictrl.currState_2_RNI2P2AZ0Z_2\
        );

    \I__3258\ : LocalMux
    port map (
            O => \N__17963\,
            I => \Lab_UT.dictrl.currState_2_RNI2P2AZ0Z_2\
        );

    \I__3257\ : LocalMux
    port map (
            O => \N__17960\,
            I => \Lab_UT.dictrl.currState_2_RNI2P2AZ0Z_2\
        );

    \I__3256\ : Odrv4
    port map (
            O => \N__17951\,
            I => \Lab_UT.dictrl.currState_2_RNI2P2AZ0Z_2\
        );

    \I__3255\ : Odrv4
    port map (
            O => \N__17946\,
            I => \Lab_UT.dictrl.currState_2_RNI2P2AZ0Z_2\
        );

    \I__3254\ : CascadeMux
    port map (
            O => \N__17929\,
            I => \N__17921\
        );

    \I__3253\ : InMux
    port map (
            O => \N__17928\,
            I => \N__17907\
        );

    \I__3252\ : InMux
    port map (
            O => \N__17927\,
            I => \N__17895\
        );

    \I__3251\ : InMux
    port map (
            O => \N__17926\,
            I => \N__17895\
        );

    \I__3250\ : InMux
    port map (
            O => \N__17925\,
            I => \N__17895\
        );

    \I__3249\ : InMux
    port map (
            O => \N__17924\,
            I => \N__17895\
        );

    \I__3248\ : InMux
    port map (
            O => \N__17921\,
            I => \N__17889\
        );

    \I__3247\ : InMux
    port map (
            O => \N__17920\,
            I => \N__17883\
        );

    \I__3246\ : InMux
    port map (
            O => \N__17919\,
            I => \N__17876\
        );

    \I__3245\ : InMux
    port map (
            O => \N__17918\,
            I => \N__17876\
        );

    \I__3244\ : InMux
    port map (
            O => \N__17917\,
            I => \N__17876\
        );

    \I__3243\ : InMux
    port map (
            O => \N__17916\,
            I => \N__17873\
        );

    \I__3242\ : InMux
    port map (
            O => \N__17915\,
            I => \N__17870\
        );

    \I__3241\ : InMux
    port map (
            O => \N__17914\,
            I => \N__17863\
        );

    \I__3240\ : InMux
    port map (
            O => \N__17913\,
            I => \N__17863\
        );

    \I__3239\ : InMux
    port map (
            O => \N__17912\,
            I => \N__17863\
        );

    \I__3238\ : InMux
    port map (
            O => \N__17911\,
            I => \N__17856\
        );

    \I__3237\ : CascadeMux
    port map (
            O => \N__17910\,
            I => \N__17851\
        );

    \I__3236\ : LocalMux
    port map (
            O => \N__17907\,
            I => \N__17848\
        );

    \I__3235\ : InMux
    port map (
            O => \N__17906\,
            I => \N__17841\
        );

    \I__3234\ : InMux
    port map (
            O => \N__17905\,
            I => \N__17841\
        );

    \I__3233\ : InMux
    port map (
            O => \N__17904\,
            I => \N__17841\
        );

    \I__3232\ : LocalMux
    port map (
            O => \N__17895\,
            I => \N__17838\
        );

    \I__3231\ : CascadeMux
    port map (
            O => \N__17894\,
            I => \N__17835\
        );

    \I__3230\ : CascadeMux
    port map (
            O => \N__17893\,
            I => \N__17832\
        );

    \I__3229\ : CascadeMux
    port map (
            O => \N__17892\,
            I => \N__17829\
        );

    \I__3228\ : LocalMux
    port map (
            O => \N__17889\,
            I => \N__17825\
        );

    \I__3227\ : InMux
    port map (
            O => \N__17888\,
            I => \N__17818\
        );

    \I__3226\ : InMux
    port map (
            O => \N__17887\,
            I => \N__17818\
        );

    \I__3225\ : InMux
    port map (
            O => \N__17886\,
            I => \N__17818\
        );

    \I__3224\ : LocalMux
    port map (
            O => \N__17883\,
            I => \N__17811\
        );

    \I__3223\ : LocalMux
    port map (
            O => \N__17876\,
            I => \N__17811\
        );

    \I__3222\ : LocalMux
    port map (
            O => \N__17873\,
            I => \N__17811\
        );

    \I__3221\ : LocalMux
    port map (
            O => \N__17870\,
            I => \N__17806\
        );

    \I__3220\ : LocalMux
    port map (
            O => \N__17863\,
            I => \N__17806\
        );

    \I__3219\ : InMux
    port map (
            O => \N__17862\,
            I => \N__17803\
        );

    \I__3218\ : InMux
    port map (
            O => \N__17861\,
            I => \N__17800\
        );

    \I__3217\ : InMux
    port map (
            O => \N__17860\,
            I => \N__17795\
        );

    \I__3216\ : InMux
    port map (
            O => \N__17859\,
            I => \N__17795\
        );

    \I__3215\ : LocalMux
    port map (
            O => \N__17856\,
            I => \N__17792\
        );

    \I__3214\ : InMux
    port map (
            O => \N__17855\,
            I => \N__17785\
        );

    \I__3213\ : InMux
    port map (
            O => \N__17854\,
            I => \N__17785\
        );

    \I__3212\ : InMux
    port map (
            O => \N__17851\,
            I => \N__17785\
        );

    \I__3211\ : Span4Mux_v
    port map (
            O => \N__17848\,
            I => \N__17778\
        );

    \I__3210\ : LocalMux
    port map (
            O => \N__17841\,
            I => \N__17778\
        );

    \I__3209\ : Span4Mux_v
    port map (
            O => \N__17838\,
            I => \N__17778\
        );

    \I__3208\ : InMux
    port map (
            O => \N__17835\,
            I => \N__17773\
        );

    \I__3207\ : InMux
    port map (
            O => \N__17832\,
            I => \N__17773\
        );

    \I__3206\ : InMux
    port map (
            O => \N__17829\,
            I => \N__17770\
        );

    \I__3205\ : InMux
    port map (
            O => \N__17828\,
            I => \N__17767\
        );

    \I__3204\ : Span4Mux_v
    port map (
            O => \N__17825\,
            I => \N__17760\
        );

    \I__3203\ : LocalMux
    port map (
            O => \N__17818\,
            I => \N__17760\
        );

    \I__3202\ : Span4Mux_v
    port map (
            O => \N__17811\,
            I => \N__17760\
        );

    \I__3201\ : Span4Mux_h
    port map (
            O => \N__17806\,
            I => \N__17753\
        );

    \I__3200\ : LocalMux
    port map (
            O => \N__17803\,
            I => \N__17753\
        );

    \I__3199\ : LocalMux
    port map (
            O => \N__17800\,
            I => \N__17753\
        );

    \I__3198\ : LocalMux
    port map (
            O => \N__17795\,
            I => \N__17750\
        );

    \I__3197\ : Span12Mux_s10_h
    port map (
            O => \N__17792\,
            I => \N__17745\
        );

    \I__3196\ : LocalMux
    port map (
            O => \N__17785\,
            I => \N__17745\
        );

    \I__3195\ : Span4Mux_h
    port map (
            O => \N__17778\,
            I => \N__17742\
        );

    \I__3194\ : LocalMux
    port map (
            O => \N__17773\,
            I => \Lab_UT_dictrl_currState_1\
        );

    \I__3193\ : LocalMux
    port map (
            O => \N__17770\,
            I => \Lab_UT_dictrl_currState_1\
        );

    \I__3192\ : LocalMux
    port map (
            O => \N__17767\,
            I => \Lab_UT_dictrl_currState_1\
        );

    \I__3191\ : Odrv4
    port map (
            O => \N__17760\,
            I => \Lab_UT_dictrl_currState_1\
        );

    \I__3190\ : Odrv4
    port map (
            O => \N__17753\,
            I => \Lab_UT_dictrl_currState_1\
        );

    \I__3189\ : Odrv4
    port map (
            O => \N__17750\,
            I => \Lab_UT_dictrl_currState_1\
        );

    \I__3188\ : Odrv12
    port map (
            O => \N__17745\,
            I => \Lab_UT_dictrl_currState_1\
        );

    \I__3187\ : Odrv4
    port map (
            O => \N__17742\,
            I => \Lab_UT_dictrl_currState_1\
        );

    \I__3186\ : InMux
    port map (
            O => \N__17725\,
            I => \N__17721\
        );

    \I__3185\ : InMux
    port map (
            O => \N__17724\,
            I => \N__17718\
        );

    \I__3184\ : LocalMux
    port map (
            O => \N__17721\,
            I => \N__17713\
        );

    \I__3183\ : LocalMux
    port map (
            O => \N__17718\,
            I => \N__17713\
        );

    \I__3182\ : Odrv12
    port map (
            O => \N__17713\,
            I => \Lab_UT.dictrl.G_19_0_a7_2\
        );

    \I__3181\ : InMux
    port map (
            O => \N__17710\,
            I => \N__17707\
        );

    \I__3180\ : LocalMux
    port map (
            O => \N__17707\,
            I => \N__17704\
        );

    \I__3179\ : Odrv4
    port map (
            O => \N__17704\,
            I => \Lab_UT.dictrl.decoder.g0_2Z0Z_2\
        );

    \I__3178\ : CascadeMux
    port map (
            O => \N__17701\,
            I => \Lab_UT_dictrl_decoder_de_cr_2_cascade_\
        );

    \I__3177\ : InMux
    port map (
            O => \N__17698\,
            I => \N__17691\
        );

    \I__3176\ : InMux
    port map (
            O => \N__17697\,
            I => \N__17688\
        );

    \I__3175\ : InMux
    port map (
            O => \N__17696\,
            I => \N__17683\
        );

    \I__3174\ : InMux
    port map (
            O => \N__17695\,
            I => \N__17683\
        );

    \I__3173\ : InMux
    port map (
            O => \N__17694\,
            I => \N__17680\
        );

    \I__3172\ : LocalMux
    port map (
            O => \N__17691\,
            I => \buart__rx_bitcount_2_rep1\
        );

    \I__3171\ : LocalMux
    port map (
            O => \N__17688\,
            I => \buart__rx_bitcount_2_rep1\
        );

    \I__3170\ : LocalMux
    port map (
            O => \N__17683\,
            I => \buart__rx_bitcount_2_rep1\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__17680\,
            I => \buart__rx_bitcount_2_rep1\
        );

    \I__3168\ : CascadeMux
    port map (
            O => \N__17671\,
            I => \Lab_UT.dictrl.decoder.g0_4_0_cascade_\
        );

    \I__3167\ : InMux
    port map (
            O => \N__17668\,
            I => \N__17664\
        );

    \I__3166\ : InMux
    port map (
            O => \N__17667\,
            I => \N__17661\
        );

    \I__3165\ : LocalMux
    port map (
            O => \N__17664\,
            I => \N__17657\
        );

    \I__3164\ : LocalMux
    port map (
            O => \N__17661\,
            I => \N__17654\
        );

    \I__3163\ : InMux
    port map (
            O => \N__17660\,
            I => \N__17651\
        );

    \I__3162\ : Span4Mux_s3_h
    port map (
            O => \N__17657\,
            I => \N__17642\
        );

    \I__3161\ : Span4Mux_s3_v
    port map (
            O => \N__17654\,
            I => \N__17642\
        );

    \I__3160\ : LocalMux
    port map (
            O => \N__17651\,
            I => \N__17642\
        );

    \I__3159\ : InMux
    port map (
            O => \N__17650\,
            I => \N__17639\
        );

    \I__3158\ : InMux
    port map (
            O => \N__17649\,
            I => \N__17636\
        );

    \I__3157\ : Odrv4
    port map (
            O => \N__17642\,
            I => \Lab_UT.dictrl.de_cr_1_0\
        );

    \I__3156\ : LocalMux
    port map (
            O => \N__17639\,
            I => \Lab_UT.dictrl.de_cr_1_0\
        );

    \I__3155\ : LocalMux
    port map (
            O => \N__17636\,
            I => \Lab_UT.dictrl.de_cr_1_0\
        );

    \I__3154\ : InMux
    port map (
            O => \N__17629\,
            I => \N__17626\
        );

    \I__3153\ : LocalMux
    port map (
            O => \N__17626\,
            I => \N__17623\
        );

    \I__3152\ : Span4Mux_h
    port map (
            O => \N__17623\,
            I => \N__17620\
        );

    \I__3151\ : Odrv4
    port map (
            O => \N__17620\,
            I => \Lab_UT.dictrl.de_cr_0\
        );

    \I__3150\ : InMux
    port map (
            O => \N__17617\,
            I => \N__17613\
        );

    \I__3149\ : InMux
    port map (
            O => \N__17616\,
            I => \N__17610\
        );

    \I__3148\ : LocalMux
    port map (
            O => \N__17613\,
            I => \N__17607\
        );

    \I__3147\ : LocalMux
    port map (
            O => \N__17610\,
            I => bu_rx_data_fast_2
        );

    \I__3146\ : Odrv4
    port map (
            O => \N__17607\,
            I => bu_rx_data_fast_2
        );

    \I__3145\ : CascadeMux
    port map (
            O => \N__17602\,
            I => \Lab_UT.dictrl.r_dicLdMtens15_1i_cascade_\
        );

    \I__3144\ : InMux
    port map (
            O => \N__17599\,
            I => \N__17596\
        );

    \I__3143\ : LocalMux
    port map (
            O => \N__17596\,
            I => \N__17593\
        );

    \I__3142\ : Span4Mux_h
    port map (
            O => \N__17593\,
            I => \N__17590\
        );

    \I__3141\ : Odrv4
    port map (
            O => \N__17590\,
            I => \Lab_UT.dictrl.currState_ret_3and\
        );

    \I__3140\ : InMux
    port map (
            O => \N__17587\,
            I => \N__17584\
        );

    \I__3139\ : LocalMux
    port map (
            O => \N__17584\,
            I => \N__17581\
        );

    \I__3138\ : Span4Mux_h
    port map (
            O => \N__17581\,
            I => \N__17578\
        );

    \I__3137\ : Span4Mux_h
    port map (
            O => \N__17578\,
            I => \N__17575\
        );

    \I__3136\ : Odrv4
    port map (
            O => \N__17575\,
            I => \Lab_UT.dictrl.currState_0_ret_28_RNOZ0Z_2\
        );

    \I__3135\ : InMux
    port map (
            O => \N__17572\,
            I => \N__17568\
        );

    \I__3134\ : InMux
    port map (
            O => \N__17571\,
            I => \N__17562\
        );

    \I__3133\ : LocalMux
    port map (
            O => \N__17568\,
            I => \N__17559\
        );

    \I__3132\ : InMux
    port map (
            O => \N__17567\,
            I => \N__17554\
        );

    \I__3131\ : InMux
    port map (
            O => \N__17566\,
            I => \N__17554\
        );

    \I__3130\ : CascadeMux
    port map (
            O => \N__17565\,
            I => \N__17549\
        );

    \I__3129\ : LocalMux
    port map (
            O => \N__17562\,
            I => \N__17543\
        );

    \I__3128\ : Span4Mux_v
    port map (
            O => \N__17559\,
            I => \N__17538\
        );

    \I__3127\ : LocalMux
    port map (
            O => \N__17554\,
            I => \N__17538\
        );

    \I__3126\ : InMux
    port map (
            O => \N__17553\,
            I => \N__17533\
        );

    \I__3125\ : InMux
    port map (
            O => \N__17552\,
            I => \N__17533\
        );

    \I__3124\ : InMux
    port map (
            O => \N__17549\,
            I => \N__17527\
        );

    \I__3123\ : InMux
    port map (
            O => \N__17548\,
            I => \N__17527\
        );

    \I__3122\ : InMux
    port map (
            O => \N__17547\,
            I => \N__17521\
        );

    \I__3121\ : InMux
    port map (
            O => \N__17546\,
            I => \N__17521\
        );

    \I__3120\ : Span4Mux_h
    port map (
            O => \N__17543\,
            I => \N__17516\
        );

    \I__3119\ : Span4Mux_h
    port map (
            O => \N__17538\,
            I => \N__17516\
        );

    \I__3118\ : LocalMux
    port map (
            O => \N__17533\,
            I => \N__17513\
        );

    \I__3117\ : InMux
    port map (
            O => \N__17532\,
            I => \N__17510\
        );

    \I__3116\ : LocalMux
    port map (
            O => \N__17527\,
            I => \N__17507\
        );

    \I__3115\ : InMux
    port map (
            O => \N__17526\,
            I => \N__17504\
        );

    \I__3114\ : LocalMux
    port map (
            O => \N__17521\,
            I => \Lab_UT.dictrl.N_8ctr\
        );

    \I__3113\ : Odrv4
    port map (
            O => \N__17516\,
            I => \Lab_UT.dictrl.N_8ctr\
        );

    \I__3112\ : Odrv4
    port map (
            O => \N__17513\,
            I => \Lab_UT.dictrl.N_8ctr\
        );

    \I__3111\ : LocalMux
    port map (
            O => \N__17510\,
            I => \Lab_UT.dictrl.N_8ctr\
        );

    \I__3110\ : Odrv12
    port map (
            O => \N__17507\,
            I => \Lab_UT.dictrl.N_8ctr\
        );

    \I__3109\ : LocalMux
    port map (
            O => \N__17504\,
            I => \Lab_UT.dictrl.N_8ctr\
        );

    \I__3108\ : CascadeMux
    port map (
            O => \N__17491\,
            I => \Lab_UT.dictrl.currState_0_ret_28_RNOZ0Z_3_cascade_\
        );

    \I__3107\ : InMux
    port map (
            O => \N__17488\,
            I => \N__17485\
        );

    \I__3106\ : LocalMux
    port map (
            O => \N__17485\,
            I => \N__17482\
        );

    \I__3105\ : Odrv4
    port map (
            O => \N__17482\,
            I => \Lab_UT.dictrl.N_8_0\
        );

    \I__3104\ : InMux
    port map (
            O => \N__17479\,
            I => \N__17476\
        );

    \I__3103\ : LocalMux
    port map (
            O => \N__17476\,
            I => \Lab_UT.dictrl.r_dicLdMtens21_1_reti\
        );

    \I__3102\ : InMux
    port map (
            O => \N__17473\,
            I => \N__17469\
        );

    \I__3101\ : InMux
    port map (
            O => \N__17472\,
            I => \N__17466\
        );

    \I__3100\ : LocalMux
    port map (
            O => \N__17469\,
            I => \N__17461\
        );

    \I__3099\ : LocalMux
    port map (
            O => \N__17466\,
            I => \N__17461\
        );

    \I__3098\ : Odrv4
    port map (
            O => \N__17461\,
            I => \Lab_UT.dictrl.decoder.de_littleA_2Z0Z_0\
        );

    \I__3097\ : CascadeMux
    port map (
            O => \N__17458\,
            I => \Lab_UT.dictrl.de_littleA_1_cascade_\
        );

    \I__3096\ : CascadeMux
    port map (
            O => \N__17455\,
            I => \Lab_UT.dictrl.N_37_0_cascade_\
        );

    \I__3095\ : InMux
    port map (
            O => \N__17452\,
            I => \N__17449\
        );

    \I__3094\ : LocalMux
    port map (
            O => \N__17449\,
            I => \N__17446\
        );

    \I__3093\ : Odrv4
    port map (
            O => \N__17446\,
            I => \Lab_UT.dictrl.g0_15_rn_1\
        );

    \I__3092\ : InMux
    port map (
            O => \N__17443\,
            I => \N__17437\
        );

    \I__3091\ : InMux
    port map (
            O => \N__17442\,
            I => \N__17437\
        );

    \I__3090\ : LocalMux
    port map (
            O => \N__17437\,
            I => \N__17434\
        );

    \I__3089\ : Span4Mux_h
    port map (
            O => \N__17434\,
            I => \N__17431\
        );

    \I__3088\ : Odrv4
    port map (
            O => \N__17431\,
            I => \Lab_UT.dictrl.G_19_0_a7_0_1\
        );

    \I__3087\ : InMux
    port map (
            O => \N__17428\,
            I => \N__17425\
        );

    \I__3086\ : LocalMux
    port map (
            O => \N__17425\,
            I => \N__17422\
        );

    \I__3085\ : Odrv12
    port map (
            O => \N__17422\,
            I => \G_19_0_a7_4_7\
        );

    \I__3084\ : InMux
    port map (
            O => \N__17419\,
            I => \N__17416\
        );

    \I__3083\ : LocalMux
    port map (
            O => \N__17416\,
            I => \N__17412\
        );

    \I__3082\ : InMux
    port map (
            O => \N__17415\,
            I => \N__17409\
        );

    \I__3081\ : Odrv4
    port map (
            O => \N__17412\,
            I => \Lab_UT.dictrl.N_17_0\
        );

    \I__3080\ : LocalMux
    port map (
            O => \N__17409\,
            I => \Lab_UT.dictrl.N_17_0\
        );

    \I__3079\ : CascadeMux
    port map (
            O => \N__17404\,
            I => \Lab_UT.dictrl.N_13_cascade_\
        );

    \I__3078\ : InMux
    port map (
            O => \N__17401\,
            I => \N__17398\
        );

    \I__3077\ : LocalMux
    port map (
            O => \N__17398\,
            I => \N__17395\
        );

    \I__3076\ : Span4Mux_v
    port map (
            O => \N__17395\,
            I => \N__17391\
        );

    \I__3075\ : InMux
    port map (
            O => \N__17394\,
            I => \N__17388\
        );

    \I__3074\ : Sp12to4
    port map (
            O => \N__17391\,
            I => \N__17383\
        );

    \I__3073\ : LocalMux
    port map (
            O => \N__17388\,
            I => \N__17383\
        );

    \I__3072\ : Span12Mux_s10_h
    port map (
            O => \N__17383\,
            I => \N__17380\
        );

    \I__3071\ : Odrv12
    port map (
            O => \N__17380\,
            I => \Lab_UT.dictrl.G_19_0_2\
        );

    \I__3070\ : CascadeMux
    port map (
            O => \N__17377\,
            I => \Lab_UT.dictrl.nextStateZ0Z_2_cascade_\
        );

    \I__3069\ : InMux
    port map (
            O => \N__17374\,
            I => \N__17371\
        );

    \I__3068\ : LocalMux
    port map (
            O => \N__17371\,
            I => \Lab_UT.dictrl.dicLdASones_rst\
        );

    \I__3067\ : CascadeMux
    port map (
            O => \N__17368\,
            I => \Lab_UT.dictrl.dicLdASones_rst_cascade_\
        );

    \I__3066\ : InMux
    port map (
            O => \N__17365\,
            I => \N__17359\
        );

    \I__3065\ : InMux
    port map (
            O => \N__17364\,
            I => \N__17359\
        );

    \I__3064\ : LocalMux
    port map (
            O => \N__17359\,
            I => \Lab_UT.dictrl.dicLdASonesZ0\
        );

    \I__3063\ : CascadeMux
    port map (
            O => \N__17356\,
            I => \N__17352\
        );

    \I__3062\ : InMux
    port map (
            O => \N__17355\,
            I => \N__17345\
        );

    \I__3061\ : InMux
    port map (
            O => \N__17352\,
            I => \N__17345\
        );

    \I__3060\ : InMux
    port map (
            O => \N__17351\,
            I => \N__17340\
        );

    \I__3059\ : InMux
    port map (
            O => \N__17350\,
            I => \N__17340\
        );

    \I__3058\ : LocalMux
    port map (
            O => \N__17345\,
            I => \Lab_UT.dictrl.N_5ctr\
        );

    \I__3057\ : LocalMux
    port map (
            O => \N__17340\,
            I => \Lab_UT.dictrl.N_5ctr\
        );

    \I__3056\ : CascadeMux
    port map (
            O => \N__17335\,
            I => \N__17332\
        );

    \I__3055\ : InMux
    port map (
            O => \N__17332\,
            I => \N__17328\
        );

    \I__3054\ : CascadeMux
    port map (
            O => \N__17331\,
            I => \N__17325\
        );

    \I__3053\ : LocalMux
    port map (
            O => \N__17328\,
            I => \N__17322\
        );

    \I__3052\ : InMux
    port map (
            O => \N__17325\,
            I => \N__17319\
        );

    \I__3051\ : Span4Mux_v
    port map (
            O => \N__17322\,
            I => \N__17316\
        );

    \I__3050\ : LocalMux
    port map (
            O => \N__17319\,
            I => \N__17313\
        );

    \I__3049\ : Odrv4
    port map (
            O => \N__17316\,
            I => \Lab_UT.dictrl.N_7ctr\
        );

    \I__3048\ : Odrv4
    port map (
            O => \N__17313\,
            I => \Lab_UT.dictrl.N_7ctr\
        );

    \I__3047\ : InMux
    port map (
            O => \N__17308\,
            I => \N__17293\
        );

    \I__3046\ : InMux
    port map (
            O => \N__17307\,
            I => \N__17293\
        );

    \I__3045\ : InMux
    port map (
            O => \N__17306\,
            I => \N__17293\
        );

    \I__3044\ : InMux
    port map (
            O => \N__17305\,
            I => \N__17293\
        );

    \I__3043\ : InMux
    port map (
            O => \N__17304\,
            I => \N__17290\
        );

    \I__3042\ : InMux
    port map (
            O => \N__17303\,
            I => \N__17285\
        );

    \I__3041\ : InMux
    port map (
            O => \N__17302\,
            I => \N__17285\
        );

    \I__3040\ : LocalMux
    port map (
            O => \N__17293\,
            I => \N__17282\
        );

    \I__3039\ : LocalMux
    port map (
            O => \N__17290\,
            I => \N__17277\
        );

    \I__3038\ : LocalMux
    port map (
            O => \N__17285\,
            I => \N__17277\
        );

    \I__3037\ : Span4Mux_v
    port map (
            O => \N__17282\,
            I => \N__17274\
        );

    \I__3036\ : Span4Mux_h
    port map (
            O => \N__17277\,
            I => \N__17271\
        );

    \I__3035\ : Odrv4
    port map (
            O => \N__17274\,
            I => \Lab_UT.dictrl.nextState_RNIGHD18Z0Z_1\
        );

    \I__3034\ : Odrv4
    port map (
            O => \N__17271\,
            I => \Lab_UT.dictrl.nextState_RNIGHD18Z0Z_1\
        );

    \I__3033\ : InMux
    port map (
            O => \N__17266\,
            I => \N__17254\
        );

    \I__3032\ : InMux
    port map (
            O => \N__17265\,
            I => \N__17247\
        );

    \I__3031\ : InMux
    port map (
            O => \N__17264\,
            I => \N__17247\
        );

    \I__3030\ : InMux
    port map (
            O => \N__17263\,
            I => \N__17247\
        );

    \I__3029\ : InMux
    port map (
            O => \N__17262\,
            I => \N__17244\
        );

    \I__3028\ : InMux
    port map (
            O => \N__17261\,
            I => \N__17241\
        );

    \I__3027\ : InMux
    port map (
            O => \N__17260\,
            I => \N__17232\
        );

    \I__3026\ : InMux
    port map (
            O => \N__17259\,
            I => \N__17232\
        );

    \I__3025\ : InMux
    port map (
            O => \N__17258\,
            I => \N__17232\
        );

    \I__3024\ : InMux
    port map (
            O => \N__17257\,
            I => \N__17232\
        );

    \I__3023\ : LocalMux
    port map (
            O => \N__17254\,
            I => \N__17225\
        );

    \I__3022\ : LocalMux
    port map (
            O => \N__17247\,
            I => \N__17225\
        );

    \I__3021\ : LocalMux
    port map (
            O => \N__17244\,
            I => \N__17222\
        );

    \I__3020\ : LocalMux
    port map (
            O => \N__17241\,
            I => \N__17216\
        );

    \I__3019\ : LocalMux
    port map (
            O => \N__17232\,
            I => \N__17216\
        );

    \I__3018\ : InMux
    port map (
            O => \N__17231\,
            I => \N__17213\
        );

    \I__3017\ : InMux
    port map (
            O => \N__17230\,
            I => \N__17210\
        );

    \I__3016\ : Span4Mux_h
    port map (
            O => \N__17225\,
            I => \N__17205\
        );

    \I__3015\ : Span4Mux_s3_h
    port map (
            O => \N__17222\,
            I => \N__17205\
        );

    \I__3014\ : InMux
    port map (
            O => \N__17221\,
            I => \N__17202\
        );

    \I__3013\ : Span4Mux_s3_h
    port map (
            O => \N__17216\,
            I => \N__17199\
        );

    \I__3012\ : LocalMux
    port map (
            O => \N__17213\,
            I => \N__17194\
        );

    \I__3011\ : LocalMux
    port map (
            O => \N__17210\,
            I => \N__17194\
        );

    \I__3010\ : Odrv4
    port map (
            O => \N__17205\,
            I => \Lab_UT.dictrl.i8_mux\
        );

    \I__3009\ : LocalMux
    port map (
            O => \N__17202\,
            I => \Lab_UT.dictrl.i8_mux\
        );

    \I__3008\ : Odrv4
    port map (
            O => \N__17199\,
            I => \Lab_UT.dictrl.i8_mux\
        );

    \I__3007\ : Odrv12
    port map (
            O => \N__17194\,
            I => \Lab_UT.dictrl.i8_mux\
        );

    \I__3006\ : CascadeMux
    port map (
            O => \N__17185\,
            I => \N__17178\
        );

    \I__3005\ : CascadeMux
    port map (
            O => \N__17184\,
            I => \N__17175\
        );

    \I__3004\ : CascadeMux
    port map (
            O => \N__17183\,
            I => \N__17172\
        );

    \I__3003\ : CascadeMux
    port map (
            O => \N__17182\,
            I => \N__17169\
        );

    \I__3002\ : CascadeMux
    port map (
            O => \N__17181\,
            I => \N__17166\
        );

    \I__3001\ : InMux
    port map (
            O => \N__17178\,
            I => \N__17161\
        );

    \I__3000\ : InMux
    port map (
            O => \N__17175\,
            I => \N__17161\
        );

    \I__2999\ : InMux
    port map (
            O => \N__17172\,
            I => \N__17156\
        );

    \I__2998\ : InMux
    port map (
            O => \N__17169\,
            I => \N__17156\
        );

    \I__2997\ : InMux
    port map (
            O => \N__17166\,
            I => \N__17153\
        );

    \I__2996\ : LocalMux
    port map (
            O => \N__17161\,
            I => \N__17148\
        );

    \I__2995\ : LocalMux
    port map (
            O => \N__17156\,
            I => \N__17148\
        );

    \I__2994\ : LocalMux
    port map (
            O => \N__17153\,
            I => \N__17145\
        );

    \I__2993\ : Span4Mux_h
    port map (
            O => \N__17148\,
            I => \N__17142\
        );

    \I__2992\ : Odrv12
    port map (
            O => \N__17145\,
            I => \Lab_UT.dictrl.currState_2_RNI1O2A_0Z0Z_1\
        );

    \I__2991\ : Odrv4
    port map (
            O => \N__17142\,
            I => \Lab_UT.dictrl.currState_2_RNI1O2A_0Z0Z_1\
        );

    \I__2990\ : InMux
    port map (
            O => \N__17137\,
            I => \N__17134\
        );

    \I__2989\ : LocalMux
    port map (
            O => \N__17134\,
            I => \N__17131\
        );

    \I__2988\ : Odrv12
    port map (
            O => \N__17131\,
            I => \Lab_UT.dictrl.g0_13_1\
        );

    \I__2987\ : InMux
    port map (
            O => \N__17128\,
            I => \N__17125\
        );

    \I__2986\ : LocalMux
    port map (
            O => \N__17125\,
            I => \Lab_UT.dictrl.g0_1\
        );

    \I__2985\ : InMux
    port map (
            O => \N__17122\,
            I => \N__17119\
        );

    \I__2984\ : LocalMux
    port map (
            O => \N__17119\,
            I => \Lab_UT.dictrl.g0_i_o4_0_0\
        );

    \I__2983\ : CascadeMux
    port map (
            O => \N__17116\,
            I => \Lab_UT.dictrl.currState_0_ret_20and_1_0_cascade_\
        );

    \I__2982\ : InMux
    port map (
            O => \N__17113\,
            I => \N__17109\
        );

    \I__2981\ : InMux
    port map (
            O => \N__17112\,
            I => \N__17106\
        );

    \I__2980\ : LocalMux
    port map (
            O => \N__17109\,
            I => \N__17103\
        );

    \I__2979\ : LocalMux
    port map (
            O => \N__17106\,
            I => \N__17100\
        );

    \I__2978\ : Span4Mux_v
    port map (
            O => \N__17103\,
            I => \N__17094\
        );

    \I__2977\ : Span4Mux_s2_h
    port map (
            O => \N__17100\,
            I => \N__17094\
        );

    \I__2976\ : InMux
    port map (
            O => \N__17099\,
            I => \N__17091\
        );

    \I__2975\ : Span4Mux_h
    port map (
            O => \N__17094\,
            I => \N__17088\
        );

    \I__2974\ : LocalMux
    port map (
            O => \N__17091\,
            I => \Lab_UT.dictrl.de_cr\
        );

    \I__2973\ : Odrv4
    port map (
            O => \N__17088\,
            I => \Lab_UT.dictrl.de_cr\
        );

    \I__2972\ : CascadeMux
    port map (
            O => \N__17083\,
            I => \N__17080\
        );

    \I__2971\ : InMux
    port map (
            O => \N__17080\,
            I => \N__17077\
        );

    \I__2970\ : LocalMux
    port map (
            O => \N__17077\,
            I => \N__17074\
        );

    \I__2969\ : Odrv4
    port map (
            O => \N__17074\,
            I => \Lab_UT.dictrl.N_13\
        );

    \I__2968\ : CascadeMux
    port map (
            O => \N__17071\,
            I => \N__17068\
        );

    \I__2967\ : InMux
    port map (
            O => \N__17068\,
            I => \N__17065\
        );

    \I__2966\ : LocalMux
    port map (
            O => \N__17065\,
            I => \N__17062\
        );

    \I__2965\ : Span4Mux_h
    port map (
            O => \N__17062\,
            I => \N__17059\
        );

    \I__2964\ : Odrv4
    port map (
            O => \N__17059\,
            I => \Lab_UT.N_91\
        );

    \I__2963\ : InMux
    port map (
            O => \N__17056\,
            I => \N__17053\
        );

    \I__2962\ : LocalMux
    port map (
            O => \N__17053\,
            I => \N__17050\
        );

    \I__2961\ : Span4Mux_h
    port map (
            O => \N__17050\,
            I => \N__17047\
        );

    \I__2960\ : Odrv4
    port map (
            O => \N__17047\,
            I => \Lab_UT.N_83\
        );

    \I__2959\ : CascadeMux
    port map (
            O => \N__17044\,
            I => \N__17034\
        );

    \I__2958\ : InMux
    port map (
            O => \N__17043\,
            I => \N__17023\
        );

    \I__2957\ : InMux
    port map (
            O => \N__17042\,
            I => \N__17023\
        );

    \I__2956\ : InMux
    port map (
            O => \N__17041\,
            I => \N__17023\
        );

    \I__2955\ : InMux
    port map (
            O => \N__17040\,
            I => \N__17023\
        );

    \I__2954\ : InMux
    port map (
            O => \N__17039\,
            I => \N__17012\
        );

    \I__2953\ : InMux
    port map (
            O => \N__17038\,
            I => \N__17012\
        );

    \I__2952\ : InMux
    port map (
            O => \N__17037\,
            I => \N__17012\
        );

    \I__2951\ : InMux
    port map (
            O => \N__17034\,
            I => \N__17012\
        );

    \I__2950\ : InMux
    port map (
            O => \N__17033\,
            I => \N__17012\
        );

    \I__2949\ : InMux
    port map (
            O => \N__17032\,
            I => \N__17009\
        );

    \I__2948\ : LocalMux
    port map (
            O => \N__17023\,
            I => \Lab_UT.Mten_at_0\
        );

    \I__2947\ : LocalMux
    port map (
            O => \N__17012\,
            I => \Lab_UT.Mten_at_0\
        );

    \I__2946\ : LocalMux
    port map (
            O => \N__17009\,
            I => \Lab_UT.Mten_at_0\
        );

    \I__2945\ : CascadeMux
    port map (
            O => \N__17002\,
            I => \N__16995\
        );

    \I__2944\ : CascadeMux
    port map (
            O => \N__17001\,
            I => \N__16991\
        );

    \I__2943\ : CascadeMux
    port map (
            O => \N__17000\,
            I => \N__16988\
        );

    \I__2942\ : CascadeMux
    port map (
            O => \N__16999\,
            I => \N__16984\
        );

    \I__2941\ : CascadeMux
    port map (
            O => \N__16998\,
            I => \N__16980\
        );

    \I__2940\ : InMux
    port map (
            O => \N__16995\,
            I => \N__16970\
        );

    \I__2939\ : InMux
    port map (
            O => \N__16994\,
            I => \N__16970\
        );

    \I__2938\ : InMux
    port map (
            O => \N__16991\,
            I => \N__16970\
        );

    \I__2937\ : InMux
    port map (
            O => \N__16988\,
            I => \N__16970\
        );

    \I__2936\ : InMux
    port map (
            O => \N__16987\,
            I => \N__16967\
        );

    \I__2935\ : InMux
    port map (
            O => \N__16984\,
            I => \N__16958\
        );

    \I__2934\ : InMux
    port map (
            O => \N__16983\,
            I => \N__16958\
        );

    \I__2933\ : InMux
    port map (
            O => \N__16980\,
            I => \N__16958\
        );

    \I__2932\ : InMux
    port map (
            O => \N__16979\,
            I => \N__16958\
        );

    \I__2931\ : LocalMux
    port map (
            O => \N__16970\,
            I => \Lab_UT.Mten_at_3\
        );

    \I__2930\ : LocalMux
    port map (
            O => \N__16967\,
            I => \Lab_UT.Mten_at_3\
        );

    \I__2929\ : LocalMux
    port map (
            O => \N__16958\,
            I => \Lab_UT.Mten_at_3\
        );

    \I__2928\ : CascadeMux
    port map (
            O => \N__16951\,
            I => \Lab_UT.Mten_at_0_cascade_\
        );

    \I__2927\ : InMux
    port map (
            O => \N__16948\,
            I => \N__16945\
        );

    \I__2926\ : LocalMux
    port map (
            O => \N__16945\,
            I => \Lab_UT.N_77\
        );

    \I__2925\ : InMux
    port map (
            O => \N__16942\,
            I => \N__16925\
        );

    \I__2924\ : InMux
    port map (
            O => \N__16941\,
            I => \N__16925\
        );

    \I__2923\ : InMux
    port map (
            O => \N__16940\,
            I => \N__16925\
        );

    \I__2922\ : InMux
    port map (
            O => \N__16939\,
            I => \N__16925\
        );

    \I__2921\ : InMux
    port map (
            O => \N__16938\,
            I => \N__16922\
        );

    \I__2920\ : InMux
    port map (
            O => \N__16937\,
            I => \N__16913\
        );

    \I__2919\ : InMux
    port map (
            O => \N__16936\,
            I => \N__16913\
        );

    \I__2918\ : InMux
    port map (
            O => \N__16935\,
            I => \N__16913\
        );

    \I__2917\ : InMux
    port map (
            O => \N__16934\,
            I => \N__16913\
        );

    \I__2916\ : LocalMux
    port map (
            O => \N__16925\,
            I => \Lab_UT.Mten_at_1\
        );

    \I__2915\ : LocalMux
    port map (
            O => \N__16922\,
            I => \Lab_UT.Mten_at_1\
        );

    \I__2914\ : LocalMux
    port map (
            O => \N__16913\,
            I => \Lab_UT.Mten_at_1\
        );

    \I__2913\ : InMux
    port map (
            O => \N__16906\,
            I => \N__16903\
        );

    \I__2912\ : LocalMux
    port map (
            O => \N__16903\,
            I => \Lab_UT.N_77_1\
        );

    \I__2911\ : InMux
    port map (
            O => \N__16900\,
            I => \N__16897\
        );

    \I__2910\ : LocalMux
    port map (
            O => \N__16897\,
            I => \uu2.bitmapZ0Z_84\
        );

    \I__2909\ : InMux
    port map (
            O => \N__16894\,
            I => \N__16891\
        );

    \I__2908\ : LocalMux
    port map (
            O => \N__16891\,
            I => \N__16888\
        );

    \I__2907\ : Span4Mux_h
    port map (
            O => \N__16888\,
            I => \N__16885\
        );

    \I__2906\ : Odrv4
    port map (
            O => \N__16885\,
            I => \Lab_UT.L3_segment4_0_i_1_5\
        );

    \I__2905\ : InMux
    port map (
            O => \N__16882\,
            I => \N__16879\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__16879\,
            I => \N__16876\
        );

    \I__2903\ : Odrv4
    port map (
            O => \N__16876\,
            I => \Lab_UT.N_65\
        );

    \I__2902\ : CascadeMux
    port map (
            O => \N__16873\,
            I => \Lab_UT.Mten_at_3_cascade_\
        );

    \I__2901\ : InMux
    port map (
            O => \N__16870\,
            I => \N__16867\
        );

    \I__2900\ : LocalMux
    port map (
            O => \N__16867\,
            I => \N__16864\
        );

    \I__2899\ : Span4Mux_h
    port map (
            O => \N__16864\,
            I => \N__16861\
        );

    \I__2898\ : Odrv4
    port map (
            O => \N__16861\,
            I => \Lab_UT.segment_1_3\
        );

    \I__2897\ : InMux
    port map (
            O => \N__16858\,
            I => \N__16852\
        );

    \I__2896\ : InMux
    port map (
            O => \N__16857\,
            I => \N__16852\
        );

    \I__2895\ : LocalMux
    port map (
            O => \N__16852\,
            I => \Lab_UT.N_69_0\
        );

    \I__2894\ : CascadeMux
    port map (
            O => \N__16849\,
            I => \Lab_UT.N_69_0_cascade_\
        );

    \I__2893\ : InMux
    port map (
            O => \N__16846\,
            I => \N__16843\
        );

    \I__2892\ : LocalMux
    port map (
            O => \N__16843\,
            I => \N__16840\
        );

    \I__2891\ : Span4Mux_h
    port map (
            O => \N__16840\,
            I => \N__16837\
        );

    \I__2890\ : Odrv4
    port map (
            O => \N__16837\,
            I => \Lab_UT.N_92\
        );

    \I__2889\ : InMux
    port map (
            O => \N__16834\,
            I => \N__16828\
        );

    \I__2888\ : InMux
    port map (
            O => \N__16833\,
            I => \N__16828\
        );

    \I__2887\ : LocalMux
    port map (
            O => \N__16828\,
            I => \Lab_UT.N_67_0\
        );

    \I__2886\ : CascadeMux
    port map (
            O => \N__16825\,
            I => \Lab_UT.N_65_2_cascade_\
        );

    \I__2885\ : InMux
    port map (
            O => \N__16822\,
            I => \N__16819\
        );

    \I__2884\ : LocalMux
    port map (
            O => \N__16819\,
            I => \Lab_UT.segment_1_2_6\
        );

    \I__2883\ : InMux
    port map (
            O => \N__16816\,
            I => \N__16813\
        );

    \I__2882\ : LocalMux
    port map (
            O => \N__16813\,
            I => \N__16810\
        );

    \I__2881\ : Odrv4
    port map (
            O => \N__16810\,
            I => \uu2.bitmapZ0Z_186\
        );

    \I__2880\ : CascadeMux
    port map (
            O => \N__16807\,
            I => \Lab_UT.N_76_2_cascade_\
        );

    \I__2879\ : InMux
    port map (
            O => \N__16804\,
            I => \N__16801\
        );

    \I__2878\ : LocalMux
    port map (
            O => \N__16801\,
            I => \uu2.bitmapZ0Z_90\
        );

    \I__2877\ : CascadeMux
    port map (
            O => \N__16798\,
            I => \N__16795\
        );

    \I__2876\ : InMux
    port map (
            O => \N__16795\,
            I => \N__16792\
        );

    \I__2875\ : LocalMux
    port map (
            O => \N__16792\,
            I => \uu2.bitmapZ0Z_218\
        );

    \I__2874\ : InMux
    port map (
            O => \N__16789\,
            I => \N__16781\
        );

    \I__2873\ : InMux
    port map (
            O => \N__16788\,
            I => \N__16781\
        );

    \I__2872\ : InMux
    port map (
            O => \N__16787\,
            I => \N__16772\
        );

    \I__2871\ : InMux
    port map (
            O => \N__16786\,
            I => \N__16772\
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__16781\,
            I => \N__16764\
        );

    \I__2869\ : InMux
    port map (
            O => \N__16780\,
            I => \N__16761\
        );

    \I__2868\ : CascadeMux
    port map (
            O => \N__16779\,
            I => \N__16758\
        );

    \I__2867\ : InMux
    port map (
            O => \N__16778\,
            I => \N__16751\
        );

    \I__2866\ : InMux
    port map (
            O => \N__16777\,
            I => \N__16751\
        );

    \I__2865\ : LocalMux
    port map (
            O => \N__16772\,
            I => \N__16748\
        );

    \I__2864\ : InMux
    port map (
            O => \N__16771\,
            I => \N__16745\
        );

    \I__2863\ : InMux
    port map (
            O => \N__16770\,
            I => \N__16740\
        );

    \I__2862\ : InMux
    port map (
            O => \N__16769\,
            I => \N__16740\
        );

    \I__2861\ : InMux
    port map (
            O => \N__16768\,
            I => \N__16737\
        );

    \I__2860\ : InMux
    port map (
            O => \N__16767\,
            I => \N__16734\
        );

    \I__2859\ : Span4Mux_h
    port map (
            O => \N__16764\,
            I => \N__16731\
        );

    \I__2858\ : LocalMux
    port map (
            O => \N__16761\,
            I => \N__16728\
        );

    \I__2857\ : InMux
    port map (
            O => \N__16758\,
            I => \N__16721\
        );

    \I__2856\ : InMux
    port map (
            O => \N__16757\,
            I => \N__16721\
        );

    \I__2855\ : InMux
    port map (
            O => \N__16756\,
            I => \N__16721\
        );

    \I__2854\ : LocalMux
    port map (
            O => \N__16751\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__2853\ : Odrv4
    port map (
            O => \N__16748\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__2852\ : LocalMux
    port map (
            O => \N__16745\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__16740\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__2850\ : LocalMux
    port map (
            O => \N__16737\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__2849\ : LocalMux
    port map (
            O => \N__16734\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__2848\ : Odrv4
    port map (
            O => \N__16731\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__2847\ : Odrv4
    port map (
            O => \N__16728\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__2846\ : LocalMux
    port map (
            O => \N__16721\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__2845\ : CascadeMux
    port map (
            O => \N__16702\,
            I => \Lab_UT.N_76_1_cascade_\
        );

    \I__2844\ : InMux
    port map (
            O => \N__16699\,
            I => \N__16696\
        );

    \I__2843\ : LocalMux
    port map (
            O => \N__16696\,
            I => \N__16693\
        );

    \I__2842\ : Span4Mux_h
    port map (
            O => \N__16693\,
            I => \N__16690\
        );

    \I__2841\ : Odrv4
    port map (
            O => \N__16690\,
            I => \uu2.bitmapZ0Z_212\
        );

    \I__2840\ : CascadeMux
    port map (
            O => \N__16687\,
            I => \Lab_UT.N_65_1_cascade_\
        );

    \I__2839\ : InMux
    port map (
            O => \N__16684\,
            I => \N__16681\
        );

    \I__2838\ : LocalMux
    port map (
            O => \N__16681\,
            I => \Lab_UT.segment_1_1_6\
        );

    \I__2837\ : InMux
    port map (
            O => \N__16678\,
            I => \N__16675\
        );

    \I__2836\ : LocalMux
    port map (
            O => \N__16675\,
            I => \uu2.bitmapZ0Z_180\
        );

    \I__2835\ : CascadeMux
    port map (
            O => \N__16672\,
            I => \Lab_UT.L3_segment2_1_2_cascade_\
        );

    \I__2834\ : CascadeMux
    port map (
            O => \N__16669\,
            I => \N__16666\
        );

    \I__2833\ : InMux
    port map (
            O => \N__16666\,
            I => \N__16663\
        );

    \I__2832\ : LocalMux
    port map (
            O => \N__16663\,
            I => \N__16660\
        );

    \I__2831\ : Span4Mux_v
    port map (
            O => \N__16660\,
            I => \N__16657\
        );

    \I__2830\ : Odrv4
    port map (
            O => \N__16657\,
            I => \uu2.bitmapZ0Z_215\
        );

    \I__2829\ : CascadeMux
    port map (
            O => \N__16654\,
            I => \Lab_UT.L3_segment2_0_i_1_0_cascade_\
        );

    \I__2828\ : InMux
    port map (
            O => \N__16651\,
            I => \N__16648\
        );

    \I__2827\ : LocalMux
    port map (
            O => \N__16648\,
            I => \uu2.bitmapZ0Z_52\
        );

    \I__2826\ : InMux
    port map (
            O => \N__16645\,
            I => \N__16636\
        );

    \I__2825\ : InMux
    port map (
            O => \N__16644\,
            I => \N__16633\
        );

    \I__2824\ : InMux
    port map (
            O => \N__16643\,
            I => \N__16628\
        );

    \I__2823\ : InMux
    port map (
            O => \N__16642\,
            I => \N__16628\
        );

    \I__2822\ : InMux
    port map (
            O => \N__16641\,
            I => \N__16622\
        );

    \I__2821\ : InMux
    port map (
            O => \N__16640\,
            I => \N__16622\
        );

    \I__2820\ : CascadeMux
    port map (
            O => \N__16639\,
            I => \N__16619\
        );

    \I__2819\ : LocalMux
    port map (
            O => \N__16636\,
            I => \N__16613\
        );

    \I__2818\ : LocalMux
    port map (
            O => \N__16633\,
            I => \N__16608\
        );

    \I__2817\ : LocalMux
    port map (
            O => \N__16628\,
            I => \N__16608\
        );

    \I__2816\ : InMux
    port map (
            O => \N__16627\,
            I => \N__16605\
        );

    \I__2815\ : LocalMux
    port map (
            O => \N__16622\,
            I => \N__16601\
        );

    \I__2814\ : InMux
    port map (
            O => \N__16619\,
            I => \N__16598\
        );

    \I__2813\ : InMux
    port map (
            O => \N__16618\,
            I => \N__16595\
        );

    \I__2812\ : InMux
    port map (
            O => \N__16617\,
            I => \N__16590\
        );

    \I__2811\ : InMux
    port map (
            O => \N__16616\,
            I => \N__16590\
        );

    \I__2810\ : Span4Mux_s3_v
    port map (
            O => \N__16613\,
            I => \N__16583\
        );

    \I__2809\ : Span4Mux_v
    port map (
            O => \N__16608\,
            I => \N__16583\
        );

    \I__2808\ : LocalMux
    port map (
            O => \N__16605\,
            I => \N__16583\
        );

    \I__2807\ : InMux
    port map (
            O => \N__16604\,
            I => \N__16580\
        );

    \I__2806\ : Span4Mux_h
    port map (
            O => \N__16601\,
            I => \N__16577\
        );

    \I__2805\ : LocalMux
    port map (
            O => \N__16598\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__2804\ : LocalMux
    port map (
            O => \N__16595\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__16590\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__2802\ : Odrv4
    port map (
            O => \N__16583\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__2801\ : LocalMux
    port map (
            O => \N__16580\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__2800\ : Odrv4
    port map (
            O => \N__16577\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__2799\ : InMux
    port map (
            O => \N__16564\,
            I => \N__16561\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__16561\,
            I => \uu2.bitmapZ0Z_308\
        );

    \I__2797\ : InMux
    port map (
            O => \N__16558\,
            I => \N__16555\
        );

    \I__2796\ : LocalMux
    port map (
            O => \N__16555\,
            I => \uu2.N_158\
        );

    \I__2795\ : CascadeMux
    port map (
            O => \N__16552\,
            I => \Lab_UT.segmentUQ_0_0_1_cascade_\
        );

    \I__2794\ : InMux
    port map (
            O => \N__16549\,
            I => \N__16546\
        );

    \I__2793\ : LocalMux
    port map (
            O => \N__16546\,
            I => \N__16540\
        );

    \I__2792\ : InMux
    port map (
            O => \N__16545\,
            I => \N__16537\
        );

    \I__2791\ : CascadeMux
    port map (
            O => \N__16544\,
            I => \N__16534\
        );

    \I__2790\ : InMux
    port map (
            O => \N__16543\,
            I => \N__16530\
        );

    \I__2789\ : Span4Mux_v
    port map (
            O => \N__16540\,
            I => \N__16525\
        );

    \I__2788\ : LocalMux
    port map (
            O => \N__16537\,
            I => \N__16525\
        );

    \I__2787\ : InMux
    port map (
            O => \N__16534\,
            I => \N__16520\
        );

    \I__2786\ : InMux
    port map (
            O => \N__16533\,
            I => \N__16520\
        );

    \I__2785\ : LocalMux
    port map (
            O => \N__16530\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__2784\ : Odrv4
    port map (
            O => \N__16525\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__16520\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__2782\ : InMux
    port map (
            O => \N__16513\,
            I => \N__16507\
        );

    \I__2781\ : InMux
    port map (
            O => \N__16512\,
            I => \N__16507\
        );

    \I__2780\ : LocalMux
    port map (
            O => \N__16507\,
            I => \N__16501\
        );

    \I__2779\ : InMux
    port map (
            O => \N__16506\,
            I => \N__16495\
        );

    \I__2778\ : InMux
    port map (
            O => \N__16505\,
            I => \N__16492\
        );

    \I__2777\ : InMux
    port map (
            O => \N__16504\,
            I => \N__16489\
        );

    \I__2776\ : Span4Mux_h
    port map (
            O => \N__16501\,
            I => \N__16486\
        );

    \I__2775\ : InMux
    port map (
            O => \N__16500\,
            I => \N__16481\
        );

    \I__2774\ : InMux
    port map (
            O => \N__16499\,
            I => \N__16481\
        );

    \I__2773\ : InMux
    port map (
            O => \N__16498\,
            I => \N__16478\
        );

    \I__2772\ : LocalMux
    port map (
            O => \N__16495\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__2771\ : LocalMux
    port map (
            O => \N__16492\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__2770\ : LocalMux
    port map (
            O => \N__16489\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__2769\ : Odrv4
    port map (
            O => \N__16486\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__2768\ : LocalMux
    port map (
            O => \N__16481\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__16478\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__2766\ : InMux
    port map (
            O => \N__16465\,
            I => \N__16462\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__16462\,
            I => \N__16458\
        );

    \I__2764\ : InMux
    port map (
            O => \N__16461\,
            I => \N__16455\
        );

    \I__2763\ : Span4Mux_v
    port map (
            O => \N__16458\,
            I => \N__16452\
        );

    \I__2762\ : LocalMux
    port map (
            O => \N__16455\,
            I => \uu2.N_41\
        );

    \I__2761\ : Odrv4
    port map (
            O => \N__16452\,
            I => \uu2.N_41\
        );

    \I__2760\ : CascadeMux
    port map (
            O => \N__16447\,
            I => \N__16443\
        );

    \I__2759\ : InMux
    port map (
            O => \N__16446\,
            I => \N__16437\
        );

    \I__2758\ : InMux
    port map (
            O => \N__16443\,
            I => \N__16434\
        );

    \I__2757\ : CascadeMux
    port map (
            O => \N__16442\,
            I => \N__16430\
        );

    \I__2756\ : InMux
    port map (
            O => \N__16441\,
            I => \N__16425\
        );

    \I__2755\ : InMux
    port map (
            O => \N__16440\,
            I => \N__16425\
        );

    \I__2754\ : LocalMux
    port map (
            O => \N__16437\,
            I => \N__16422\
        );

    \I__2753\ : LocalMux
    port map (
            O => \N__16434\,
            I => \N__16419\
        );

    \I__2752\ : InMux
    port map (
            O => \N__16433\,
            I => \N__16416\
        );

    \I__2751\ : InMux
    port map (
            O => \N__16430\,
            I => \N__16413\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__16425\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__2749\ : Odrv4
    port map (
            O => \N__16422\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__2748\ : Odrv4
    port map (
            O => \N__16419\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__16416\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__2746\ : LocalMux
    port map (
            O => \N__16413\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__2745\ : CascadeMux
    port map (
            O => \N__16402\,
            I => \uu2.N_41_cascade_\
        );

    \I__2744\ : InMux
    port map (
            O => \N__16399\,
            I => \N__16392\
        );

    \I__2743\ : InMux
    port map (
            O => \N__16398\,
            I => \N__16392\
        );

    \I__2742\ : CascadeMux
    port map (
            O => \N__16397\,
            I => \N__16389\
        );

    \I__2741\ : LocalMux
    port map (
            O => \N__16392\,
            I => \N__16385\
        );

    \I__2740\ : InMux
    port map (
            O => \N__16389\,
            I => \N__16380\
        );

    \I__2739\ : InMux
    port map (
            O => \N__16388\,
            I => \N__16380\
        );

    \I__2738\ : Odrv4
    port map (
            O => \N__16385\,
            I => \uu2.N_43\
        );

    \I__2737\ : LocalMux
    port map (
            O => \N__16380\,
            I => \uu2.N_43\
        );

    \I__2736\ : InMux
    port map (
            O => \N__16375\,
            I => \N__16371\
        );

    \I__2735\ : CascadeMux
    port map (
            O => \N__16374\,
            I => \N__16368\
        );

    \I__2734\ : LocalMux
    port map (
            O => \N__16371\,
            I => \N__16365\
        );

    \I__2733\ : InMux
    port map (
            O => \N__16368\,
            I => \N__16358\
        );

    \I__2732\ : Span4Mux_v
    port map (
            O => \N__16365\,
            I => \N__16355\
        );

    \I__2731\ : InMux
    port map (
            O => \N__16364\,
            I => \N__16346\
        );

    \I__2730\ : InMux
    port map (
            O => \N__16363\,
            I => \N__16346\
        );

    \I__2729\ : InMux
    port map (
            O => \N__16362\,
            I => \N__16346\
        );

    \I__2728\ : InMux
    port map (
            O => \N__16361\,
            I => \N__16346\
        );

    \I__2727\ : LocalMux
    port map (
            O => \N__16358\,
            I => \uu2.N_40\
        );

    \I__2726\ : Odrv4
    port map (
            O => \N__16355\,
            I => \uu2.N_40\
        );

    \I__2725\ : LocalMux
    port map (
            O => \N__16346\,
            I => \uu2.N_40\
        );

    \I__2724\ : CascadeMux
    port map (
            O => \N__16339\,
            I => \uu2.N_43_cascade_\
        );

    \I__2723\ : CascadeMux
    port map (
            O => \N__16336\,
            I => \N__16333\
        );

    \I__2722\ : InMux
    port map (
            O => \N__16333\,
            I => \N__16326\
        );

    \I__2721\ : InMux
    port map (
            O => \N__16332\,
            I => \N__16323\
        );

    \I__2720\ : InMux
    port map (
            O => \N__16331\,
            I => \N__16316\
        );

    \I__2719\ : InMux
    port map (
            O => \N__16330\,
            I => \N__16316\
        );

    \I__2718\ : InMux
    port map (
            O => \N__16329\,
            I => \N__16316\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__16326\,
            I => \N__16311\
        );

    \I__2716\ : LocalMux
    port map (
            O => \N__16323\,
            I => \N__16311\
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__16316\,
            I => \uu2.w_addr_displaying_RNIFCPV4Z0Z_8\
        );

    \I__2714\ : Odrv4
    port map (
            O => \N__16311\,
            I => \uu2.w_addr_displaying_RNIFCPV4Z0Z_8\
        );

    \I__2713\ : CascadeMux
    port map (
            O => \N__16306\,
            I => \uu2.w_addr_displaying_RNIFCPV4Z0Z_8_cascade_\
        );

    \I__2712\ : CEMux
    port map (
            O => \N__16303\,
            I => \N__16300\
        );

    \I__2711\ : LocalMux
    port map (
            O => \N__16300\,
            I => \N__16297\
        );

    \I__2710\ : Odrv4
    port map (
            O => \N__16297\,
            I => \uu2.N_36_0\
        );

    \I__2709\ : InMux
    port map (
            O => \N__16294\,
            I => \N__16291\
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__16291\,
            I => \Lab_UT.L3_segment2_1_1\
        );

    \I__2707\ : CascadeMux
    port map (
            O => \N__16288\,
            I => \Lab_UT.L3_segment2_0_i_1_3_cascade_\
        );

    \I__2706\ : CascadeMux
    port map (
            O => \N__16285\,
            I => \uu2.un3_w_addr_user_4_cascade_\
        );

    \I__2705\ : InMux
    port map (
            O => \N__16282\,
            I => \N__16279\
        );

    \I__2704\ : LocalMux
    port map (
            O => \N__16279\,
            I => \uu2.un3_w_addr_user_5\
        );

    \I__2703\ : InMux
    port map (
            O => \N__16276\,
            I => \N__16268\
        );

    \I__2702\ : InMux
    port map (
            O => \N__16275\,
            I => \N__16260\
        );

    \I__2701\ : InMux
    port map (
            O => \N__16274\,
            I => \N__16260\
        );

    \I__2700\ : InMux
    port map (
            O => \N__16273\,
            I => \N__16260\
        );

    \I__2699\ : CascadeMux
    port map (
            O => \N__16272\,
            I => \N__16247\
        );

    \I__2698\ : InMux
    port map (
            O => \N__16271\,
            I => \N__16244\
        );

    \I__2697\ : LocalMux
    port map (
            O => \N__16268\,
            I => \N__16241\
        );

    \I__2696\ : InMux
    port map (
            O => \N__16267\,
            I => \N__16238\
        );

    \I__2695\ : LocalMux
    port map (
            O => \N__16260\,
            I => \N__16235\
        );

    \I__2694\ : InMux
    port map (
            O => \N__16259\,
            I => \N__16232\
        );

    \I__2693\ : InMux
    port map (
            O => \N__16258\,
            I => \N__16227\
        );

    \I__2692\ : InMux
    port map (
            O => \N__16257\,
            I => \N__16227\
        );

    \I__2691\ : InMux
    port map (
            O => \N__16256\,
            I => \N__16218\
        );

    \I__2690\ : InMux
    port map (
            O => \N__16255\,
            I => \N__16218\
        );

    \I__2689\ : InMux
    port map (
            O => \N__16254\,
            I => \N__16218\
        );

    \I__2688\ : InMux
    port map (
            O => \N__16253\,
            I => \N__16218\
        );

    \I__2687\ : InMux
    port map (
            O => \N__16252\,
            I => \N__16209\
        );

    \I__2686\ : InMux
    port map (
            O => \N__16251\,
            I => \N__16209\
        );

    \I__2685\ : InMux
    port map (
            O => \N__16250\,
            I => \N__16209\
        );

    \I__2684\ : InMux
    port map (
            O => \N__16247\,
            I => \N__16209\
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__16244\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__2682\ : Odrv4
    port map (
            O => \N__16241\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__16238\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__2680\ : Odrv4
    port map (
            O => \N__16235\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__16232\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__2678\ : LocalMux
    port map (
            O => \N__16227\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__16218\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__2676\ : LocalMux
    port map (
            O => \N__16209\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__2675\ : CascadeMux
    port map (
            O => \N__16192\,
            I => \N__16189\
        );

    \I__2674\ : InMux
    port map (
            O => \N__16189\,
            I => \N__16186\
        );

    \I__2673\ : LocalMux
    port map (
            O => \N__16186\,
            I => \N__16183\
        );

    \I__2672\ : Odrv12
    port map (
            O => \N__16183\,
            I => \uu2.mem0.w_addr_3\
        );

    \I__2671\ : CascadeMux
    port map (
            O => \N__16180\,
            I => \uu2.vbuf_w_addr_user.un448_ci_0_cascade_\
        );

    \I__2670\ : InMux
    port map (
            O => \N__16177\,
            I => \N__16174\
        );

    \I__2669\ : LocalMux
    port map (
            O => \N__16174\,
            I => \N__16169\
        );

    \I__2668\ : InMux
    port map (
            O => \N__16173\,
            I => \N__16164\
        );

    \I__2667\ : InMux
    port map (
            O => \N__16172\,
            I => \N__16164\
        );

    \I__2666\ : Odrv4
    port map (
            O => \N__16169\,
            I => \uu2.w_addr_userZ0Z_8\
        );

    \I__2665\ : LocalMux
    port map (
            O => \N__16164\,
            I => \uu2.w_addr_userZ0Z_8\
        );

    \I__2664\ : InMux
    port map (
            O => \N__16159\,
            I => \N__16156\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__16156\,
            I => \N__16152\
        );

    \I__2662\ : CascadeMux
    port map (
            O => \N__16155\,
            I => \N__16147\
        );

    \I__2661\ : Span4Mux_h
    port map (
            O => \N__16152\,
            I => \N__16144\
        );

    \I__2660\ : InMux
    port map (
            O => \N__16151\,
            I => \N__16137\
        );

    \I__2659\ : InMux
    port map (
            O => \N__16150\,
            I => \N__16137\
        );

    \I__2658\ : InMux
    port map (
            O => \N__16147\,
            I => \N__16137\
        );

    \I__2657\ : Odrv4
    port map (
            O => \N__16144\,
            I => \uu2.w_addr_userZ0Z_7\
        );

    \I__2656\ : LocalMux
    port map (
            O => \N__16137\,
            I => \uu2.w_addr_userZ0Z_7\
        );

    \I__2655\ : InMux
    port map (
            O => \N__16132\,
            I => \N__16122\
        );

    \I__2654\ : InMux
    port map (
            O => \N__16131\,
            I => \N__16122\
        );

    \I__2653\ : InMux
    port map (
            O => \N__16130\,
            I => \N__16122\
        );

    \I__2652\ : InMux
    port map (
            O => \N__16129\,
            I => \N__16115\
        );

    \I__2651\ : LocalMux
    port map (
            O => \N__16122\,
            I => \N__16112\
        );

    \I__2650\ : CascadeMux
    port map (
            O => \N__16121\,
            I => \N__16105\
        );

    \I__2649\ : InMux
    port map (
            O => \N__16120\,
            I => \N__16098\
        );

    \I__2648\ : InMux
    port map (
            O => \N__16119\,
            I => \N__16098\
        );

    \I__2647\ : InMux
    port map (
            O => \N__16118\,
            I => \N__16095\
        );

    \I__2646\ : LocalMux
    port map (
            O => \N__16115\,
            I => \N__16092\
        );

    \I__2645\ : Span4Mux_h
    port map (
            O => \N__16112\,
            I => \N__16089\
        );

    \I__2644\ : InMux
    port map (
            O => \N__16111\,
            I => \N__16084\
        );

    \I__2643\ : InMux
    port map (
            O => \N__16110\,
            I => \N__16084\
        );

    \I__2642\ : InMux
    port map (
            O => \N__16109\,
            I => \N__16081\
        );

    \I__2641\ : InMux
    port map (
            O => \N__16108\,
            I => \N__16072\
        );

    \I__2640\ : InMux
    port map (
            O => \N__16105\,
            I => \N__16072\
        );

    \I__2639\ : InMux
    port map (
            O => \N__16104\,
            I => \N__16072\
        );

    \I__2638\ : InMux
    port map (
            O => \N__16103\,
            I => \N__16072\
        );

    \I__2637\ : LocalMux
    port map (
            O => \N__16098\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__16095\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__2635\ : Odrv4
    port map (
            O => \N__16092\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__2634\ : Odrv4
    port map (
            O => \N__16089\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__16084\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__2632\ : LocalMux
    port map (
            O => \N__16081\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__2631\ : LocalMux
    port map (
            O => \N__16072\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__2630\ : CascadeMux
    port map (
            O => \N__16057\,
            I => \N__16054\
        );

    \I__2629\ : InMux
    port map (
            O => \N__16054\,
            I => \N__16047\
        );

    \I__2628\ : InMux
    port map (
            O => \N__16053\,
            I => \N__16047\
        );

    \I__2627\ : CascadeMux
    port map (
            O => \N__16052\,
            I => \N__16044\
        );

    \I__2626\ : LocalMux
    port map (
            O => \N__16047\,
            I => \N__16041\
        );

    \I__2625\ : InMux
    port map (
            O => \N__16044\,
            I => \N__16038\
        );

    \I__2624\ : Odrv4
    port map (
            O => \N__16041\,
            I => \uu2.N_39\
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__16038\,
            I => \uu2.N_39\
        );

    \I__2622\ : InMux
    port map (
            O => \N__16033\,
            I => \N__16030\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__16030\,
            I => \N__16026\
        );

    \I__2620\ : InMux
    port map (
            O => \N__16029\,
            I => \N__16023\
        );

    \I__2619\ : Span4Mux_h
    port map (
            O => \N__16026\,
            I => \N__16020\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__16023\,
            I => \Lab_UT.uu0.l_countZ0Z_13\
        );

    \I__2617\ : Odrv4
    port map (
            O => \N__16020\,
            I => \Lab_UT.uu0.l_countZ0Z_13\
        );

    \I__2616\ : CascadeMux
    port map (
            O => \N__16015\,
            I => \Lab_UT.uu0.un143_ci_0_cascade_\
        );

    \I__2615\ : CascadeMux
    port map (
            O => \N__16012\,
            I => \Lab_UT.uu0.un154_ci_9_cascade_\
        );

    \I__2614\ : InMux
    port map (
            O => \N__16009\,
            I => \N__16006\
        );

    \I__2613\ : LocalMux
    port map (
            O => \N__16006\,
            I => \N__16001\
        );

    \I__2612\ : InMux
    port map (
            O => \N__16005\,
            I => \N__15996\
        );

    \I__2611\ : InMux
    port map (
            O => \N__16004\,
            I => \N__15996\
        );

    \I__2610\ : Span4Mux_h
    port map (
            O => \N__16001\,
            I => \N__15993\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__15996\,
            I => \Lab_UT.uu0.l_countZ0Z_12\
        );

    \I__2608\ : Odrv4
    port map (
            O => \N__15993\,
            I => \Lab_UT.uu0.l_countZ0Z_12\
        );

    \I__2607\ : CascadeMux
    port map (
            O => \N__15988\,
            I => \N__15985\
        );

    \I__2606\ : InMux
    port map (
            O => \N__15985\,
            I => \N__15982\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__15982\,
            I => \Lab_UT.uu0.un165_ci_0\
        );

    \I__2604\ : InMux
    port map (
            O => \N__15979\,
            I => \N__15955\
        );

    \I__2603\ : InMux
    port map (
            O => \N__15978\,
            I => \N__15955\
        );

    \I__2602\ : InMux
    port map (
            O => \N__15977\,
            I => \N__15955\
        );

    \I__2601\ : InMux
    port map (
            O => \N__15976\,
            I => \N__15955\
        );

    \I__2600\ : InMux
    port map (
            O => \N__15975\,
            I => \N__15955\
        );

    \I__2599\ : InMux
    port map (
            O => \N__15974\,
            I => \N__15955\
        );

    \I__2598\ : InMux
    port map (
            O => \N__15973\,
            I => \N__15955\
        );

    \I__2597\ : InMux
    port map (
            O => \N__15972\,
            I => \N__15955\
        );

    \I__2596\ : LocalMux
    port map (
            O => \N__15955\,
            I => \N__15951\
        );

    \I__2595\ : InMux
    port map (
            O => \N__15954\,
            I => \N__15948\
        );

    \I__2594\ : Odrv4
    port map (
            O => \N__15951\,
            I => \buart.Z_rx.N_27_0_i\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__15948\,
            I => \buart.Z_rx.N_27_0_i\
        );

    \I__2592\ : CascadeMux
    port map (
            O => \N__15943\,
            I => \N__15938\
        );

    \I__2591\ : CascadeMux
    port map (
            O => \N__15942\,
            I => \N__15935\
        );

    \I__2590\ : CascadeMux
    port map (
            O => \N__15941\,
            I => \N__15932\
        );

    \I__2589\ : InMux
    port map (
            O => \N__15938\,
            I => \N__15902\
        );

    \I__2588\ : InMux
    port map (
            O => \N__15935\,
            I => \N__15902\
        );

    \I__2587\ : InMux
    port map (
            O => \N__15932\,
            I => \N__15902\
        );

    \I__2586\ : InMux
    port map (
            O => \N__15931\,
            I => \N__15902\
        );

    \I__2585\ : InMux
    port map (
            O => \N__15930\,
            I => \N__15902\
        );

    \I__2584\ : InMux
    port map (
            O => \N__15929\,
            I => \N__15902\
        );

    \I__2583\ : InMux
    port map (
            O => \N__15928\,
            I => \N__15902\
        );

    \I__2582\ : InMux
    port map (
            O => \N__15927\,
            I => \N__15902\
        );

    \I__2581\ : InMux
    port map (
            O => \N__15926\,
            I => \N__15897\
        );

    \I__2580\ : InMux
    port map (
            O => \N__15925\,
            I => \N__15897\
        );

    \I__2579\ : InMux
    port map (
            O => \N__15924\,
            I => \N__15892\
        );

    \I__2578\ : InMux
    port map (
            O => \N__15923\,
            I => \N__15892\
        );

    \I__2577\ : InMux
    port map (
            O => \N__15922\,
            I => \N__15887\
        );

    \I__2576\ : InMux
    port map (
            O => \N__15921\,
            I => \N__15887\
        );

    \I__2575\ : InMux
    port map (
            O => \N__15920\,
            I => \N__15882\
        );

    \I__2574\ : InMux
    port map (
            O => \N__15919\,
            I => \N__15882\
        );

    \I__2573\ : LocalMux
    port map (
            O => \N__15902\,
            I => \buart.Z_rx.startbit\
        );

    \I__2572\ : LocalMux
    port map (
            O => \N__15897\,
            I => \buart.Z_rx.startbit\
        );

    \I__2571\ : LocalMux
    port map (
            O => \N__15892\,
            I => \buart.Z_rx.startbit\
        );

    \I__2570\ : LocalMux
    port map (
            O => \N__15887\,
            I => \buart.Z_rx.startbit\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__15882\,
            I => \buart.Z_rx.startbit\
        );

    \I__2568\ : CEMux
    port map (
            O => \N__15871\,
            I => \N__15867\
        );

    \I__2567\ : CEMux
    port map (
            O => \N__15870\,
            I => \N__15864\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__15867\,
            I => \N__15861\
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__15864\,
            I => \N__15858\
        );

    \I__2564\ : Span4Mux_h
    port map (
            O => \N__15861\,
            I => \N__15855\
        );

    \I__2563\ : Span4Mux_h
    port map (
            O => \N__15858\,
            I => \N__15852\
        );

    \I__2562\ : Span4Mux_s1_v
    port map (
            O => \N__15855\,
            I => \N__15849\
        );

    \I__2561\ : Odrv4
    port map (
            O => \N__15852\,
            I => \buart.Z_rx.bitcounte_0_0\
        );

    \I__2560\ : Odrv4
    port map (
            O => \N__15849\,
            I => \buart.Z_rx.bitcounte_0_0\
        );

    \I__2559\ : InMux
    port map (
            O => \N__15844\,
            I => \N__15839\
        );

    \I__2558\ : CascadeMux
    port map (
            O => \N__15843\,
            I => \N__15832\
        );

    \I__2557\ : InMux
    port map (
            O => \N__15842\,
            I => \N__15829\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__15839\,
            I => \N__15826\
        );

    \I__2555\ : InMux
    port map (
            O => \N__15838\,
            I => \N__15817\
        );

    \I__2554\ : InMux
    port map (
            O => \N__15837\,
            I => \N__15817\
        );

    \I__2553\ : InMux
    port map (
            O => \N__15836\,
            I => \N__15817\
        );

    \I__2552\ : InMux
    port map (
            O => \N__15835\,
            I => \N__15817\
        );

    \I__2551\ : InMux
    port map (
            O => \N__15832\,
            I => \N__15814\
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__15829\,
            I => \buart__rx_bitcount_0\
        );

    \I__2549\ : Odrv4
    port map (
            O => \N__15826\,
            I => \buart__rx_bitcount_0\
        );

    \I__2548\ : LocalMux
    port map (
            O => \N__15817\,
            I => \buart__rx_bitcount_0\
        );

    \I__2547\ : LocalMux
    port map (
            O => \N__15814\,
            I => \buart__rx_bitcount_0\
        );

    \I__2546\ : InMux
    port map (
            O => \N__15805\,
            I => \N__15800\
        );

    \I__2545\ : CascadeMux
    port map (
            O => \N__15804\,
            I => \N__15797\
        );

    \I__2544\ : InMux
    port map (
            O => \N__15803\,
            I => \N__15790\
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__15800\,
            I => \N__15787\
        );

    \I__2542\ : InMux
    port map (
            O => \N__15797\,
            I => \N__15784\
        );

    \I__2541\ : InMux
    port map (
            O => \N__15796\,
            I => \N__15781\
        );

    \I__2540\ : InMux
    port map (
            O => \N__15795\,
            I => \N__15778\
        );

    \I__2539\ : InMux
    port map (
            O => \N__15794\,
            I => \N__15773\
        );

    \I__2538\ : InMux
    port map (
            O => \N__15793\,
            I => \N__15773\
        );

    \I__2537\ : LocalMux
    port map (
            O => \N__15790\,
            I => \buart__rx_bitcount_1\
        );

    \I__2536\ : Odrv4
    port map (
            O => \N__15787\,
            I => \buart__rx_bitcount_1\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__15784\,
            I => \buart__rx_bitcount_1\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__15781\,
            I => \buart__rx_bitcount_1\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__15778\,
            I => \buart__rx_bitcount_1\
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__15773\,
            I => \buart__rx_bitcount_1\
        );

    \I__2531\ : CascadeMux
    port map (
            O => \N__15760\,
            I => \N__15757\
        );

    \I__2530\ : InMux
    port map (
            O => \N__15757\,
            I => \N__15754\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__15754\,
            I => \N__15751\
        );

    \I__2528\ : Odrv4
    port map (
            O => \N__15751\,
            I => \buart.Z_rx.bitcount_cry_0_THRU_CO\
        );

    \I__2527\ : InMux
    port map (
            O => \N__15748\,
            I => \buart.Z_rx.bitcount_cry_0\
        );

    \I__2526\ : CascadeMux
    port map (
            O => \N__15745\,
            I => \N__15741\
        );

    \I__2525\ : CascadeMux
    port map (
            O => \N__15744\,
            I => \N__15737\
        );

    \I__2524\ : InMux
    port map (
            O => \N__15741\,
            I => \N__15730\
        );

    \I__2523\ : InMux
    port map (
            O => \N__15740\,
            I => \N__15730\
        );

    \I__2522\ : InMux
    port map (
            O => \N__15737\,
            I => \N__15730\
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__15730\,
            I => \N__15727\
        );

    \I__2520\ : Odrv4
    port map (
            O => \N__15727\,
            I => \buart.Z_rx.bitcount_cry_1_THRU_CO\
        );

    \I__2519\ : InMux
    port map (
            O => \N__15724\,
            I => \buart.Z_rx.bitcount_cry_1\
        );

    \I__2518\ : CascadeMux
    port map (
            O => \N__15721\,
            I => \N__15717\
        );

    \I__2517\ : InMux
    port map (
            O => \N__15720\,
            I => \N__15712\
        );

    \I__2516\ : InMux
    port map (
            O => \N__15717\,
            I => \N__15712\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__15712\,
            I => \N__15709\
        );

    \I__2514\ : Odrv4
    port map (
            O => \N__15709\,
            I => \buart.Z_rx.bitcount_cry_2_THRU_CO\
        );

    \I__2513\ : InMux
    port map (
            O => \N__15706\,
            I => \buart.Z_rx.bitcount_cry_2\
        );

    \I__2512\ : InMux
    port map (
            O => \N__15703\,
            I => \buart.Z_rx.bitcount_cry_3\
        );

    \I__2511\ : CascadeMux
    port map (
            O => \N__15700\,
            I => \N__15696\
        );

    \I__2510\ : InMux
    port map (
            O => \N__15699\,
            I => \N__15691\
        );

    \I__2509\ : InMux
    port map (
            O => \N__15696\,
            I => \N__15691\
        );

    \I__2508\ : LocalMux
    port map (
            O => \N__15691\,
            I => \N__15688\
        );

    \I__2507\ : Odrv12
    port map (
            O => \N__15688\,
            I => \buart.Z_rx.bitcount_cry_3_THRU_CO\
        );

    \I__2506\ : CascadeMux
    port map (
            O => \N__15685\,
            I => \N__15682\
        );

    \I__2505\ : InMux
    port map (
            O => \N__15682\,
            I => \N__15676\
        );

    \I__2504\ : InMux
    port map (
            O => \N__15681\,
            I => \N__15676\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__15676\,
            I => \buart__rx_bitcount_fast_4\
        );

    \I__2502\ : InMux
    port map (
            O => \N__15673\,
            I => \N__15670\
        );

    \I__2501\ : LocalMux
    port map (
            O => \N__15670\,
            I => \N__15666\
        );

    \I__2500\ : InMux
    port map (
            O => \N__15669\,
            I => \N__15663\
        );

    \I__2499\ : Odrv4
    port map (
            O => \N__15666\,
            I => \buart__rx_bitcount_fast_3\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__15663\,
            I => \buart__rx_bitcount_fast_3\
        );

    \I__2497\ : InMux
    port map (
            O => \N__15658\,
            I => \N__15655\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__15655\,
            I => \Lab_UT.dictrl.decoder.g0_6_1\
        );

    \I__2495\ : CascadeMux
    port map (
            O => \N__15652\,
            I => \buart.Z_rx.un1_sample_0_cascade_\
        );

    \I__2494\ : IoInMux
    port map (
            O => \N__15649\,
            I => \N__15646\
        );

    \I__2493\ : LocalMux
    port map (
            O => \N__15646\,
            I => \N__15643\
        );

    \I__2492\ : Odrv4
    port map (
            O => \N__15643\,
            I => \buart.Z_rx.sample\
        );

    \I__2491\ : CascadeMux
    port map (
            O => \N__15640\,
            I => \buart.Z_rx.idle_0_cascade_\
        );

    \I__2490\ : InMux
    port map (
            O => \N__15637\,
            I => \N__15633\
        );

    \I__2489\ : InMux
    port map (
            O => \N__15636\,
            I => \N__15630\
        );

    \I__2488\ : LocalMux
    port map (
            O => \N__15633\,
            I => \buart.Z_rx.idle\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__15630\,
            I => \buart.Z_rx.idle\
        );

    \I__2486\ : CascadeMux
    port map (
            O => \N__15625\,
            I => \N__15621\
        );

    \I__2485\ : InMux
    port map (
            O => \N__15624\,
            I => \N__15616\
        );

    \I__2484\ : InMux
    port map (
            O => \N__15621\,
            I => \N__15613\
        );

    \I__2483\ : InMux
    port map (
            O => \N__15620\,
            I => \N__15608\
        );

    \I__2482\ : InMux
    port map (
            O => \N__15619\,
            I => \N__15608\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__15616\,
            I => \buart.Z_rx.ser_clk\
        );

    \I__2480\ : LocalMux
    port map (
            O => \N__15613\,
            I => \buart.Z_rx.ser_clk\
        );

    \I__2479\ : LocalMux
    port map (
            O => \N__15608\,
            I => \buart.Z_rx.ser_clk\
        );

    \I__2478\ : CascadeMux
    port map (
            O => \N__15601\,
            I => \buart.Z_rx.idle_cascade_\
        );

    \I__2477\ : CascadeMux
    port map (
            O => \N__15598\,
            I => \Lab_UT_dictrl_decoder_de_cr_1_cascade_\
        );

    \I__2476\ : InMux
    port map (
            O => \N__15595\,
            I => \N__15592\
        );

    \I__2475\ : LocalMux
    port map (
            O => \N__15592\,
            I => \Lab_UT.dictrl.N_30\
        );

    \I__2474\ : InMux
    port map (
            O => \N__15589\,
            I => \N__15586\
        );

    \I__2473\ : LocalMux
    port map (
            O => \N__15586\,
            I => \Lab_UT.dictrl.N_41_mux\
        );

    \I__2472\ : CascadeMux
    port map (
            O => \N__15583\,
            I => \N__15579\
        );

    \I__2471\ : InMux
    port map (
            O => \N__15582\,
            I => \N__15576\
        );

    \I__2470\ : InMux
    port map (
            O => \N__15579\,
            I => \N__15572\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__15576\,
            I => \N__15569\
        );

    \I__2468\ : CascadeMux
    port map (
            O => \N__15575\,
            I => \N__15565\
        );

    \I__2467\ : LocalMux
    port map (
            O => \N__15572\,
            I => \N__15562\
        );

    \I__2466\ : Span4Mux_h
    port map (
            O => \N__15569\,
            I => \N__15559\
        );

    \I__2465\ : InMux
    port map (
            O => \N__15568\,
            I => \N__15554\
        );

    \I__2464\ : InMux
    port map (
            O => \N__15565\,
            I => \N__15554\
        );

    \I__2463\ : Span4Mux_h
    port map (
            O => \N__15562\,
            I => \N__15551\
        );

    \I__2462\ : Odrv4
    port map (
            O => \N__15559\,
            I => \Lab_UT.dictrl.N_34\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__15554\,
            I => \Lab_UT.dictrl.N_34\
        );

    \I__2460\ : Odrv4
    port map (
            O => \N__15551\,
            I => \Lab_UT.dictrl.N_34\
        );

    \I__2459\ : CascadeMux
    port map (
            O => \N__15544\,
            I => \Lab_UT.dictrl.N_31_cascade_\
        );

    \I__2458\ : InMux
    port map (
            O => \N__15541\,
            I => \N__15538\
        );

    \I__2457\ : LocalMux
    port map (
            O => \N__15538\,
            I => \N__15534\
        );

    \I__2456\ : InMux
    port map (
            O => \N__15537\,
            I => \N__15531\
        );

    \I__2455\ : Span4Mux_s2_h
    port map (
            O => \N__15534\,
            I => \N__15528\
        );

    \I__2454\ : LocalMux
    port map (
            O => \N__15531\,
            I => \N__15525\
        );

    \I__2453\ : Span4Mux_v
    port map (
            O => \N__15528\,
            I => \N__15522\
        );

    \I__2452\ : Odrv12
    port map (
            O => \N__15525\,
            I => \Lab_UT.dictrl.nextState_0_2\
        );

    \I__2451\ : Odrv4
    port map (
            O => \N__15522\,
            I => \Lab_UT.dictrl.nextState_0_2\
        );

    \I__2450\ : CEMux
    port map (
            O => \N__15517\,
            I => \N__15514\
        );

    \I__2449\ : LocalMux
    port map (
            O => \N__15514\,
            I => \N__15510\
        );

    \I__2448\ : CEMux
    port map (
            O => \N__15513\,
            I => \N__15507\
        );

    \I__2447\ : Span4Mux_v
    port map (
            O => \N__15510\,
            I => \N__15504\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__15507\,
            I => \N__15501\
        );

    \I__2445\ : Odrv4
    port map (
            O => \N__15504\,
            I => \Lab_UT.dictrl.currState_0_ret_29_RNIDFRSEEZ0\
        );

    \I__2444\ : Odrv12
    port map (
            O => \N__15501\,
            I => \Lab_UT.dictrl.currState_0_ret_29_RNIDFRSEEZ0\
        );

    \I__2443\ : CascadeMux
    port map (
            O => \N__15496\,
            I => \N__15493\
        );

    \I__2442\ : InMux
    port map (
            O => \N__15493\,
            I => \N__15490\
        );

    \I__2441\ : LocalMux
    port map (
            O => \N__15490\,
            I => \buart__rx_bitcount_fast_2\
        );

    \I__2440\ : CascadeMux
    port map (
            O => \N__15487\,
            I => \Lab_UT.dictrl.r_dicLdMtens20_0_cascade_\
        );

    \I__2439\ : InMux
    port map (
            O => \N__15484\,
            I => \N__15477\
        );

    \I__2438\ : InMux
    port map (
            O => \N__15483\,
            I => \N__15467\
        );

    \I__2437\ : InMux
    port map (
            O => \N__15482\,
            I => \N__15467\
        );

    \I__2436\ : InMux
    port map (
            O => \N__15481\,
            I => \N__15462\
        );

    \I__2435\ : InMux
    port map (
            O => \N__15480\,
            I => \N__15462\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__15477\,
            I => \N__15459\
        );

    \I__2433\ : InMux
    port map (
            O => \N__15476\,
            I => \N__15456\
        );

    \I__2432\ : InMux
    port map (
            O => \N__15475\,
            I => \N__15451\
        );

    \I__2431\ : InMux
    port map (
            O => \N__15474\,
            I => \N__15451\
        );

    \I__2430\ : InMux
    port map (
            O => \N__15473\,
            I => \N__15446\
        );

    \I__2429\ : InMux
    port map (
            O => \N__15472\,
            I => \N__15446\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__15467\,
            I => \N__15443\
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__15462\,
            I => \N__15440\
        );

    \I__2426\ : Span4Mux_h
    port map (
            O => \N__15459\,
            I => \N__15435\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__15456\,
            I => \N__15435\
        );

    \I__2424\ : LocalMux
    port map (
            O => \N__15451\,
            I => \N__15429\
        );

    \I__2423\ : LocalMux
    port map (
            O => \N__15446\,
            I => \N__15429\
        );

    \I__2422\ : Span4Mux_s3_h
    port map (
            O => \N__15443\,
            I => \N__15424\
        );

    \I__2421\ : Span4Mux_h
    port map (
            O => \N__15440\,
            I => \N__15424\
        );

    \I__2420\ : Span4Mux_h
    port map (
            O => \N__15435\,
            I => \N__15421\
        );

    \I__2419\ : InMux
    port map (
            O => \N__15434\,
            I => \N__15418\
        );

    \I__2418\ : Odrv12
    port map (
            O => \N__15429\,
            I => \Lab_UT.dictrl.N_6ctr\
        );

    \I__2417\ : Odrv4
    port map (
            O => \N__15424\,
            I => \Lab_UT.dictrl.N_6ctr\
        );

    \I__2416\ : Odrv4
    port map (
            O => \N__15421\,
            I => \Lab_UT.dictrl.N_6ctr\
        );

    \I__2415\ : LocalMux
    port map (
            O => \N__15418\,
            I => \Lab_UT.dictrl.N_6ctr\
        );

    \I__2414\ : InMux
    port map (
            O => \N__15409\,
            I => \N__15406\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__15406\,
            I => \Lab_UT.dictrl.r_dicLdMtens22_2_reti\
        );

    \I__2412\ : InMux
    port map (
            O => \N__15403\,
            I => \N__15400\
        );

    \I__2411\ : LocalMux
    port map (
            O => \N__15400\,
            I => \N__15397\
        );

    \I__2410\ : Odrv12
    port map (
            O => \N__15397\,
            I => \Lab_UT.dictrl.N_7_1_0\
        );

    \I__2409\ : CascadeMux
    port map (
            O => \N__15394\,
            I => \Lab_UT.dictrl.r_dicLdMtens22_2_reti_cascade_\
        );

    \I__2408\ : InMux
    port map (
            O => \N__15391\,
            I => \N__15388\
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__15388\,
            I => \Lab_UT.dictrl.g0_0_3\
        );

    \I__2406\ : InMux
    port map (
            O => \N__15385\,
            I => \N__15381\
        );

    \I__2405\ : InMux
    port map (
            O => \N__15384\,
            I => \N__15378\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__15381\,
            I => \N__15374\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__15378\,
            I => \N__15371\
        );

    \I__2402\ : InMux
    port map (
            O => \N__15377\,
            I => \N__15368\
        );

    \I__2401\ : Span4Mux_h
    port map (
            O => \N__15374\,
            I => \N__15363\
        );

    \I__2400\ : Span4Mux_v
    port map (
            O => \N__15371\,
            I => \N__15363\
        );

    \I__2399\ : LocalMux
    port map (
            O => \N__15368\,
            I => \Lab_UT.dictrl.N_10ctr\
        );

    \I__2398\ : Odrv4
    port map (
            O => \N__15363\,
            I => \Lab_UT.dictrl.N_10ctr\
        );

    \I__2397\ : InMux
    port map (
            O => \N__15358\,
            I => \N__15352\
        );

    \I__2396\ : InMux
    port map (
            O => \N__15357\,
            I => \N__15352\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__15352\,
            I => \Lab_UT.dictrl.r_dicLdMtens22_4_0\
        );

    \I__2394\ : InMux
    port map (
            O => \N__15349\,
            I => \N__15346\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__15346\,
            I => \N__15343\
        );

    \I__2392\ : Span4Mux_h
    port map (
            O => \N__15343\,
            I => \N__15340\
        );

    \I__2391\ : Odrv4
    port map (
            O => \N__15340\,
            I => \N_7\
        );

    \I__2390\ : CascadeMux
    port map (
            O => \N__15337\,
            I => \N__15333\
        );

    \I__2389\ : InMux
    port map (
            O => \N__15336\,
            I => \N__15330\
        );

    \I__2388\ : InMux
    port map (
            O => \N__15333\,
            I => \N__15327\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__15330\,
            I => \N__15324\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__15327\,
            I => \N__15321\
        );

    \I__2385\ : Span4Mux_s3_h
    port map (
            O => \N__15324\,
            I => \N__15317\
        );

    \I__2384\ : Span4Mux_h
    port map (
            O => \N__15321\,
            I => \N__15314\
        );

    \I__2383\ : InMux
    port map (
            O => \N__15320\,
            I => \N__15311\
        );

    \I__2382\ : Odrv4
    port map (
            O => \N__15317\,
            I => \Lab_UT.dictrl.N_20\
        );

    \I__2381\ : Odrv4
    port map (
            O => \N__15314\,
            I => \Lab_UT.dictrl.N_20\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__15311\,
            I => \Lab_UT.dictrl.N_20\
        );

    \I__2379\ : InMux
    port map (
            O => \N__15304\,
            I => \N__15301\
        );

    \I__2378\ : LocalMux
    port map (
            O => \N__15301\,
            I => \N__15298\
        );

    \I__2377\ : Span4Mux_h
    port map (
            O => \N__15298\,
            I => \N__15294\
        );

    \I__2376\ : InMux
    port map (
            O => \N__15297\,
            I => \N__15291\
        );

    \I__2375\ : Odrv4
    port map (
            O => \N__15294\,
            I => \Lab_UT.dictrl.de_littleA\
        );

    \I__2374\ : LocalMux
    port map (
            O => \N__15291\,
            I => \Lab_UT.dictrl.de_littleA\
        );

    \I__2373\ : CascadeMux
    port map (
            O => \N__15286\,
            I => \Lab_UT.dictrl.g2_cascade_\
        );

    \I__2372\ : CascadeMux
    port map (
            O => \N__15283\,
            I => \Lab_UT.dictrl.nextState_RNO_9Z0Z_1_cascade_\
        );

    \I__2371\ : InMux
    port map (
            O => \N__15280\,
            I => \N__15276\
        );

    \I__2370\ : InMux
    port map (
            O => \N__15279\,
            I => \N__15273\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__15276\,
            I => \N__15268\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__15273\,
            I => \N__15268\
        );

    \I__2367\ : Span4Mux_v
    port map (
            O => \N__15268\,
            I => \N__15265\
        );

    \I__2366\ : Odrv4
    port map (
            O => \N__15265\,
            I => \Lab_UT.dictrl.g0_i_a4_1\
        );

    \I__2365\ : CascadeMux
    port map (
            O => \N__15262\,
            I => \Lab_UT.dictrl.nextState_RNO_4Z0Z_1_cascade_\
        );

    \I__2364\ : InMux
    port map (
            O => \N__15259\,
            I => \N__15256\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__15256\,
            I => \Lab_UT.dictrl.nextState_RNO_3Z0Z_1\
        );

    \I__2362\ : InMux
    port map (
            O => \N__15253\,
            I => \N__15250\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__15250\,
            I => \N__15247\
        );

    \I__2360\ : Odrv12
    port map (
            O => \N__15247\,
            I => \Lab_UT.dictrl.g0_i_o4_5\
        );

    \I__2359\ : InMux
    port map (
            O => \N__15244\,
            I => \N__15241\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__15241\,
            I => \Lab_UT.dictrl.N_11\
        );

    \I__2357\ : InMux
    port map (
            O => \N__15238\,
            I => \N__15235\
        );

    \I__2356\ : LocalMux
    port map (
            O => \N__15235\,
            I => \Lab_UT.dictrl.N_18_0\
        );

    \I__2355\ : CascadeMux
    port map (
            O => \N__15232\,
            I => \N__15229\
        );

    \I__2354\ : InMux
    port map (
            O => \N__15229\,
            I => \N__15226\
        );

    \I__2353\ : LocalMux
    port map (
            O => \N__15226\,
            I => \Lab_UT.dictrl.g1_3_0\
        );

    \I__2352\ : InMux
    port map (
            O => \N__15223\,
            I => \N__15220\
        );

    \I__2351\ : LocalMux
    port map (
            O => \N__15220\,
            I => \N__15217\
        );

    \I__2350\ : Odrv4
    port map (
            O => \N__15217\,
            I => \Lab_UT.dictrl.N_13_0\
        );

    \I__2349\ : CascadeMux
    port map (
            O => \N__15214\,
            I => \Lab_UT.dictrl.g1_4_0_cascade_\
        );

    \I__2348\ : InMux
    port map (
            O => \N__15211\,
            I => \N__15208\
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__15208\,
            I => \Lab_UT.dictrl.N_14\
        );

    \I__2346\ : CascadeMux
    port map (
            O => \N__15205\,
            I => \Lab_UT.dictrl.N_36_0_cascade_\
        );

    \I__2345\ : CascadeMux
    port map (
            O => \N__15202\,
            I => \Lab_UT.dictrl.nextStateZ0Z_3_cascade_\
        );

    \I__2344\ : InMux
    port map (
            O => \N__15199\,
            I => \N__15196\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__15196\,
            I => \Lab_UT.dictrl.r_dicLdMtens21_1\
        );

    \I__2342\ : InMux
    port map (
            O => \N__15193\,
            I => \N__15189\
        );

    \I__2341\ : InMux
    port map (
            O => \N__15192\,
            I => \N__15186\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__15189\,
            I => \Lab_UT.dictrl.N_18\
        );

    \I__2339\ : LocalMux
    port map (
            O => \N__15186\,
            I => \Lab_UT.dictrl.N_18\
        );

    \I__2338\ : InMux
    port map (
            O => \N__15181\,
            I => \N__15178\
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__15178\,
            I => \Lab_UT.dictrl.N_33\
        );

    \I__2336\ : InMux
    port map (
            O => \N__15175\,
            I => \N__15172\
        );

    \I__2335\ : LocalMux
    port map (
            O => \N__15172\,
            I => \Lab_UT.dictrl.N_1607_0_0\
        );

    \I__2334\ : InMux
    port map (
            O => \N__15169\,
            I => \N__15166\
        );

    \I__2333\ : LocalMux
    port map (
            O => \N__15166\,
            I => \Lab_UT.dictrl.N_10_0_0\
        );

    \I__2332\ : InMux
    port map (
            O => \N__15163\,
            I => \N__15160\
        );

    \I__2331\ : LocalMux
    port map (
            O => \N__15160\,
            I => \Lab_UT.dictrl.g1\
        );

    \I__2330\ : CascadeMux
    port map (
            O => \N__15157\,
            I => \N__15154\
        );

    \I__2329\ : InMux
    port map (
            O => \N__15154\,
            I => \N__15151\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__15151\,
            I => \N__15148\
        );

    \I__2327\ : Span4Mux_h
    port map (
            O => \N__15148\,
            I => \N__15145\
        );

    \I__2326\ : Odrv4
    port map (
            O => \N__15145\,
            I => \Lab_UT.dictrl.N_1614_0\
        );

    \I__2325\ : CascadeMux
    port map (
            O => \N__15142\,
            I => \N__15139\
        );

    \I__2324\ : InMux
    port map (
            O => \N__15139\,
            I => \N__15136\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__15136\,
            I => \Lab_UT.dictrl.N_26\
        );

    \I__2322\ : InMux
    port map (
            O => \N__15133\,
            I => \N__15130\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__15130\,
            I => \Lab_UT.dictrl.un1_currState_6\
        );

    \I__2320\ : InMux
    port map (
            O => \N__15127\,
            I => \N__15121\
        );

    \I__2319\ : InMux
    port map (
            O => \N__15126\,
            I => \N__15121\
        );

    \I__2318\ : LocalMux
    port map (
            O => \N__15121\,
            I => \Lab_UT.dictrl.r_enableZ0Z1\
        );

    \I__2317\ : InMux
    port map (
            O => \N__15118\,
            I => \N__15112\
        );

    \I__2316\ : InMux
    port map (
            O => \N__15117\,
            I => \N__15112\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__15112\,
            I => \N__15104\
        );

    \I__2314\ : InMux
    port map (
            O => \N__15111\,
            I => \N__15099\
        );

    \I__2313\ : InMux
    port map (
            O => \N__15110\,
            I => \N__15099\
        );

    \I__2312\ : InMux
    port map (
            O => \N__15109\,
            I => \N__15096\
        );

    \I__2311\ : InMux
    port map (
            O => \N__15108\,
            I => \N__15091\
        );

    \I__2310\ : InMux
    port map (
            O => \N__15107\,
            I => \N__15091\
        );

    \I__2309\ : Sp12to4
    port map (
            O => \N__15104\,
            I => \N__15088\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__15099\,
            I => \N__15081\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__15096\,
            I => \N__15081\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__15091\,
            I => \N__15081\
        );

    \I__2305\ : Odrv12
    port map (
            O => \N__15088\,
            I => \Lab_UT.dictrl.enableSeg3\
        );

    \I__2304\ : Odrv4
    port map (
            O => \N__15081\,
            I => \Lab_UT.dictrl.enableSeg3\
        );

    \I__2303\ : CascadeMux
    port map (
            O => \N__15076\,
            I => \N__15073\
        );

    \I__2302\ : InMux
    port map (
            O => \N__15073\,
            I => \N__15067\
        );

    \I__2301\ : InMux
    port map (
            O => \N__15072\,
            I => \N__15067\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__15067\,
            I => \Lab_UT.dictrl.r_enableZ0Z3\
        );

    \I__2299\ : CascadeMux
    port map (
            O => \N__15064\,
            I => \N__15061\
        );

    \I__2298\ : InMux
    port map (
            O => \N__15061\,
            I => \N__15056\
        );

    \I__2297\ : InMux
    port map (
            O => \N__15060\,
            I => \N__15050\
        );

    \I__2296\ : InMux
    port map (
            O => \N__15059\,
            I => \N__15050\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__15056\,
            I => \N__15047\
        );

    \I__2294\ : InMux
    port map (
            O => \N__15055\,
            I => \N__15044\
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__15050\,
            I => \N__15041\
        );

    \I__2292\ : Span4Mux_v
    port map (
            O => \N__15047\,
            I => \N__15035\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__15044\,
            I => \N__15032\
        );

    \I__2290\ : Span4Mux_h
    port map (
            O => \N__15041\,
            I => \N__15029\
        );

    \I__2289\ : InMux
    port map (
            O => \N__15040\,
            I => \N__15022\
        );

    \I__2288\ : InMux
    port map (
            O => \N__15039\,
            I => \N__15022\
        );

    \I__2287\ : InMux
    port map (
            O => \N__15038\,
            I => \N__15022\
        );

    \I__2286\ : Odrv4
    port map (
            O => \N__15035\,
            I => \Lab_UT.dictrl.enableSeg4\
        );

    \I__2285\ : Odrv4
    port map (
            O => \N__15032\,
            I => \Lab_UT.dictrl.enableSeg4\
        );

    \I__2284\ : Odrv4
    port map (
            O => \N__15029\,
            I => \Lab_UT.dictrl.enableSeg4\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__15022\,
            I => \Lab_UT.dictrl.enableSeg4\
        );

    \I__2282\ : InMux
    port map (
            O => \N__15013\,
            I => \N__15010\
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__15010\,
            I => \N__15007\
        );

    \I__2280\ : Odrv4
    port map (
            O => \N__15007\,
            I => \Lab_UT.dictrl.un1_currState_7\
        );

    \I__2279\ : CascadeMux
    port map (
            O => \N__15004\,
            I => \N__15001\
        );

    \I__2278\ : InMux
    port map (
            O => \N__15001\,
            I => \N__14995\
        );

    \I__2277\ : InMux
    port map (
            O => \N__15000\,
            I => \N__14995\
        );

    \I__2276\ : LocalMux
    port map (
            O => \N__14995\,
            I => \Lab_UT.dictrl.r_enableZ0Z4\
        );

    \I__2275\ : InMux
    port map (
            O => \N__14992\,
            I => \N__14989\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__14989\,
            I => \N__14986\
        );

    \I__2273\ : Odrv4
    port map (
            O => \N__14986\,
            I => \Lab_UT.dictrl.N_1605_1_0\
        );

    \I__2272\ : CascadeMux
    port map (
            O => \N__14983\,
            I => \Lab_UT.N_76_cascade_\
        );

    \I__2271\ : CascadeMux
    port map (
            O => \N__14980\,
            I => \N__14977\
        );

    \I__2270\ : InMux
    port map (
            O => \N__14977\,
            I => \N__14974\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__14974\,
            I => \N__14971\
        );

    \I__2268\ : Odrv4
    port map (
            O => \N__14971\,
            I => \uu2.bitmapZ0Z_194\
        );

    \I__2267\ : CascadeMux
    port map (
            O => \N__14968\,
            I => \Lab_UT.L3_segment4_1_1_cascade_\
        );

    \I__2266\ : InMux
    port map (
            O => \N__14965\,
            I => \N__14962\
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__14962\,
            I => \N__14959\
        );

    \I__2264\ : Odrv4
    port map (
            O => \N__14959\,
            I => \uu2.bitmapZ0Z_69\
        );

    \I__2263\ : InMux
    port map (
            O => \N__14956\,
            I => \N__14953\
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__14953\,
            I => \Lab_UT.L3_segment4_1_0\
        );

    \I__2261\ : InMux
    port map (
            O => \N__14950\,
            I => \N__14947\
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__14947\,
            I => \N__14944\
        );

    \I__2259\ : Odrv4
    port map (
            O => \N__14944\,
            I => \uu2.bitmapZ0Z_34\
        );

    \I__2258\ : CascadeMux
    port map (
            O => \N__14941\,
            I => \Lab_UT.segment_1_6_cascade_\
        );

    \I__2257\ : InMux
    port map (
            O => \N__14938\,
            I => \N__14935\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__14935\,
            I => \N__14932\
        );

    \I__2255\ : Odrv12
    port map (
            O => \N__14932\,
            I => \uu2.bitmapZ0Z_162\
        );

    \I__2254\ : InMux
    port map (
            O => \N__14929\,
            I => \N__14926\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__14926\,
            I => \N__14923\
        );

    \I__2252\ : Odrv4
    port map (
            O => \N__14923\,
            I => \uu2.bitmap_pmux_sn_N_15\
        );

    \I__2251\ : InMux
    port map (
            O => \N__14920\,
            I => \N__14910\
        );

    \I__2250\ : InMux
    port map (
            O => \N__14919\,
            I => \N__14910\
        );

    \I__2249\ : InMux
    port map (
            O => \N__14918\,
            I => \N__14910\
        );

    \I__2248\ : InMux
    port map (
            O => \N__14917\,
            I => \N__14903\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__14910\,
            I => \N__14900\
        );

    \I__2246\ : InMux
    port map (
            O => \N__14909\,
            I => \N__14891\
        );

    \I__2245\ : InMux
    port map (
            O => \N__14908\,
            I => \N__14891\
        );

    \I__2244\ : InMux
    port map (
            O => \N__14907\,
            I => \N__14891\
        );

    \I__2243\ : InMux
    port map (
            O => \N__14906\,
            I => \N__14888\
        );

    \I__2242\ : LocalMux
    port map (
            O => \N__14903\,
            I => \N__14885\
        );

    \I__2241\ : Span4Mux_h
    port map (
            O => \N__14900\,
            I => \N__14882\
        );

    \I__2240\ : InMux
    port map (
            O => \N__14899\,
            I => \N__14877\
        );

    \I__2239\ : InMux
    port map (
            O => \N__14898\,
            I => \N__14877\
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__14891\,
            I => \N__14874\
        );

    \I__2237\ : LocalMux
    port map (
            O => \N__14888\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__2236\ : Odrv12
    port map (
            O => \N__14885\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__2235\ : Odrv4
    port map (
            O => \N__14882\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__14877\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__2233\ : Odrv4
    port map (
            O => \N__14874\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__2232\ : InMux
    port map (
            O => \N__14863\,
            I => \N__14860\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__14860\,
            I => \N__14857\
        );

    \I__2230\ : Odrv4
    port map (
            O => \N__14857\,
            I => \Lab_UT.L3_segment3_0_i_1_0\
        );

    \I__2229\ : InMux
    port map (
            O => \N__14854\,
            I => \N__14851\
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__14851\,
            I => \N__14848\
        );

    \I__2227\ : Odrv4
    port map (
            O => \N__14848\,
            I => \Lab_UT.L3_segment3_0_i_1_3\
        );

    \I__2226\ : CascadeMux
    port map (
            O => \N__14845\,
            I => \Lab_UT.L3_segment3_1_2_cascade_\
        );

    \I__2225\ : InMux
    port map (
            O => \N__14842\,
            I => \N__14826\
        );

    \I__2224\ : InMux
    port map (
            O => \N__14841\,
            I => \N__14826\
        );

    \I__2223\ : InMux
    port map (
            O => \N__14840\,
            I => \N__14826\
        );

    \I__2222\ : InMux
    port map (
            O => \N__14839\,
            I => \N__14826\
        );

    \I__2221\ : InMux
    port map (
            O => \N__14838\,
            I => \N__14817\
        );

    \I__2220\ : InMux
    port map (
            O => \N__14837\,
            I => \N__14817\
        );

    \I__2219\ : InMux
    port map (
            O => \N__14836\,
            I => \N__14817\
        );

    \I__2218\ : InMux
    port map (
            O => \N__14835\,
            I => \N__14817\
        );

    \I__2217\ : LocalMux
    port map (
            O => \N__14826\,
            I => \Lab_UT.Mone_at_0\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__14817\,
            I => \Lab_UT.Mone_at_0\
        );

    \I__2215\ : CascadeMux
    port map (
            O => \N__14812\,
            I => \N__14805\
        );

    \I__2214\ : CascadeMux
    port map (
            O => \N__14811\,
            I => \N__14800\
        );

    \I__2213\ : CascadeMux
    port map (
            O => \N__14810\,
            I => \N__14797\
        );

    \I__2212\ : InMux
    port map (
            O => \N__14809\,
            I => \N__14786\
        );

    \I__2211\ : InMux
    port map (
            O => \N__14808\,
            I => \N__14786\
        );

    \I__2210\ : InMux
    port map (
            O => \N__14805\,
            I => \N__14786\
        );

    \I__2209\ : InMux
    port map (
            O => \N__14804\,
            I => \N__14786\
        );

    \I__2208\ : InMux
    port map (
            O => \N__14803\,
            I => \N__14777\
        );

    \I__2207\ : InMux
    port map (
            O => \N__14800\,
            I => \N__14777\
        );

    \I__2206\ : InMux
    port map (
            O => \N__14797\,
            I => \N__14777\
        );

    \I__2205\ : InMux
    port map (
            O => \N__14796\,
            I => \N__14777\
        );

    \I__2204\ : InMux
    port map (
            O => \N__14795\,
            I => \N__14774\
        );

    \I__2203\ : LocalMux
    port map (
            O => \N__14786\,
            I => \Lab_UT.Mone_at_3\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__14777\,
            I => \Lab_UT.Mone_at_3\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__14774\,
            I => \Lab_UT.Mone_at_3\
        );

    \I__2200\ : CascadeMux
    port map (
            O => \N__14767\,
            I => \N__14758\
        );

    \I__2199\ : CascadeMux
    port map (
            O => \N__14766\,
            I => \N__14755\
        );

    \I__2198\ : CascadeMux
    port map (
            O => \N__14765\,
            I => \N__14751\
        );

    \I__2197\ : InMux
    port map (
            O => \N__14764\,
            I => \N__14742\
        );

    \I__2196\ : InMux
    port map (
            O => \N__14763\,
            I => \N__14742\
        );

    \I__2195\ : InMux
    port map (
            O => \N__14762\,
            I => \N__14742\
        );

    \I__2194\ : InMux
    port map (
            O => \N__14761\,
            I => \N__14742\
        );

    \I__2193\ : InMux
    port map (
            O => \N__14758\,
            I => \N__14733\
        );

    \I__2192\ : InMux
    port map (
            O => \N__14755\,
            I => \N__14733\
        );

    \I__2191\ : InMux
    port map (
            O => \N__14754\,
            I => \N__14733\
        );

    \I__2190\ : InMux
    port map (
            O => \N__14751\,
            I => \N__14733\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__14742\,
            I => \Lab_UT.Mone_at_2\
        );

    \I__2188\ : LocalMux
    port map (
            O => \N__14733\,
            I => \Lab_UT.Mone_at_2\
        );

    \I__2187\ : CascadeMux
    port map (
            O => \N__14728\,
            I => \N__14724\
        );

    \I__2186\ : CascadeMux
    port map (
            O => \N__14727\,
            I => \N__14721\
        );

    \I__2185\ : InMux
    port map (
            O => \N__14724\,
            I => \N__14706\
        );

    \I__2184\ : InMux
    port map (
            O => \N__14721\,
            I => \N__14706\
        );

    \I__2183\ : InMux
    port map (
            O => \N__14720\,
            I => \N__14706\
        );

    \I__2182\ : InMux
    port map (
            O => \N__14719\,
            I => \N__14706\
        );

    \I__2181\ : InMux
    port map (
            O => \N__14718\,
            I => \N__14697\
        );

    \I__2180\ : InMux
    port map (
            O => \N__14717\,
            I => \N__14697\
        );

    \I__2179\ : InMux
    port map (
            O => \N__14716\,
            I => \N__14697\
        );

    \I__2178\ : InMux
    port map (
            O => \N__14715\,
            I => \N__14697\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__14706\,
            I => \Lab_UT.Mone_at_1\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__14697\,
            I => \Lab_UT.Mone_at_1\
        );

    \I__2175\ : CascadeMux
    port map (
            O => \N__14692\,
            I => \Lab_UT.L3_segment3_1_1_cascade_\
        );

    \I__2174\ : InMux
    port map (
            O => \N__14689\,
            I => \N__14686\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__14686\,
            I => \uu2.bitmapZ0Z_203\
        );

    \I__2172\ : InMux
    port map (
            O => \N__14683\,
            I => \N__14680\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__14680\,
            I => \uu2.bitmapZ0Z_75\
        );

    \I__2170\ : InMux
    port map (
            O => \N__14677\,
            I => \N__14674\
        );

    \I__2169\ : LocalMux
    port map (
            O => \N__14674\,
            I => \uu2.bitmap_pmux_24_bm_1\
        );

    \I__2168\ : InMux
    port map (
            O => \N__14671\,
            I => \N__14668\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__14668\,
            I => \N__14665\
        );

    \I__2166\ : Span4Mux_v
    port map (
            O => \N__14665\,
            I => \N__14662\
        );

    \I__2165\ : Odrv4
    port map (
            O => \N__14662\,
            I => \uu2.N_48\
        );

    \I__2164\ : InMux
    port map (
            O => \N__14659\,
            I => \N__14656\
        );

    \I__2163\ : LocalMux
    port map (
            O => \N__14656\,
            I => \uu2.bitmap_pmux_24_am_1\
        );

    \I__2162\ : InMux
    port map (
            O => \N__14653\,
            I => \N__14650\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__14650\,
            I => \uu2.bitmapZ0Z_87\
        );

    \I__2160\ : CascadeMux
    port map (
            O => \N__14647\,
            I => \uu2.N_386_cascade_\
        );

    \I__2159\ : CascadeMux
    port map (
            O => \N__14644\,
            I => \uu2.w_addr_displaying_nesr_RNI1JET2Z0Z_7_cascade_\
        );

    \I__2158\ : InMux
    port map (
            O => \N__14641\,
            I => \N__14635\
        );

    \I__2157\ : InMux
    port map (
            O => \N__14640\,
            I => \N__14635\
        );

    \I__2156\ : LocalMux
    port map (
            O => \N__14635\,
            I => \uu2.bitmapZ0Z_314\
        );

    \I__2155\ : InMux
    port map (
            O => \N__14632\,
            I => \N__14629\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__14629\,
            I => \uu2.bitmap_pmux_23_ns_1\
        );

    \I__2153\ : InMux
    port map (
            O => \N__14626\,
            I => \N__14623\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__14623\,
            I => \uu2.bitmap_pmux_sn_N_20\
        );

    \I__2151\ : InMux
    port map (
            O => \N__14620\,
            I => \N__14617\
        );

    \I__2150\ : LocalMux
    port map (
            O => \N__14617\,
            I => \N__14614\
        );

    \I__2149\ : Odrv4
    port map (
            O => \N__14614\,
            I => \uu2.bitmapZ0Z_168\
        );

    \I__2148\ : CascadeMux
    port map (
            O => \N__14611\,
            I => \uu2.N_17_cascade_\
        );

    \I__2147\ : InMux
    port map (
            O => \N__14608\,
            I => \N__14605\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__14605\,
            I => \uu2.bitmap_RNIELSJ2Z0Z_111\
        );

    \I__2145\ : InMux
    port map (
            O => \N__14602\,
            I => \N__14599\
        );

    \I__2144\ : LocalMux
    port map (
            O => \N__14599\,
            I => \uu2.bitmap_pmux_sn_N_54_mux\
        );

    \I__2143\ : InMux
    port map (
            O => \N__14596\,
            I => \N__14593\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__14593\,
            I => \uu2.bitmapZ0Z_111\
        );

    \I__2141\ : CascadeMux
    port map (
            O => \N__14590\,
            I => \N__14586\
        );

    \I__2140\ : InMux
    port map (
            O => \N__14589\,
            I => \N__14578\
        );

    \I__2139\ : InMux
    port map (
            O => \N__14586\,
            I => \N__14578\
        );

    \I__2138\ : InMux
    port map (
            O => \N__14585\,
            I => \N__14578\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__14578\,
            I => \N__14575\
        );

    \I__2136\ : Span4Mux_v
    port map (
            O => \N__14575\,
            I => \N__14572\
        );

    \I__2135\ : Odrv4
    port map (
            O => \N__14572\,
            I => \uu2.bitmap_pmux_sn_N_33\
        );

    \I__2134\ : CascadeMux
    port map (
            O => \N__14569\,
            I => \uu2.N_39_cascade_\
        );

    \I__2133\ : CascadeMux
    port map (
            O => \N__14566\,
            I => \resetGen.reset_count_2_0_4_cascade_\
        );

    \I__2132\ : CascadeMux
    port map (
            O => \N__14563\,
            I => \N__14560\
        );

    \I__2131\ : InMux
    port map (
            O => \N__14560\,
            I => \N__14557\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__14557\,
            I => \N__14554\
        );

    \I__2129\ : Odrv4
    port map (
            O => \N__14554\,
            I => \uu2.mem0.w_addr_2\
        );

    \I__2128\ : CascadeMux
    port map (
            O => \N__14551\,
            I => \N__14548\
        );

    \I__2127\ : InMux
    port map (
            O => \N__14548\,
            I => \N__14545\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__14545\,
            I => \N__14542\
        );

    \I__2125\ : Span4Mux_s3_h
    port map (
            O => \N__14542\,
            I => \N__14539\
        );

    \I__2124\ : Odrv4
    port map (
            O => \N__14539\,
            I => \uu2.mem0.w_addr_4\
        );

    \I__2123\ : CascadeMux
    port map (
            O => \N__14536\,
            I => \N__14533\
        );

    \I__2122\ : InMux
    port map (
            O => \N__14533\,
            I => \N__14530\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__14530\,
            I => \N__14527\
        );

    \I__2120\ : Odrv4
    port map (
            O => \N__14527\,
            I => \uu2.mem0.w_addr_5\
        );

    \I__2119\ : CascadeMux
    port map (
            O => \N__14524\,
            I => \N__14521\
        );

    \I__2118\ : InMux
    port map (
            O => \N__14521\,
            I => \N__14518\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__14518\,
            I => \N__14515\
        );

    \I__2116\ : Odrv12
    port map (
            O => \N__14515\,
            I => \uu2.mem0.w_addr_6\
        );

    \I__2115\ : CascadeMux
    port map (
            O => \N__14512\,
            I => \Lab_UT.dictrl.decoder.g0Z0Z_7_cascade_\
        );

    \I__2114\ : InMux
    port map (
            O => \N__14509\,
            I => \N__14505\
        );

    \I__2113\ : CascadeMux
    port map (
            O => \N__14508\,
            I => \N__14502\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__14505\,
            I => \N__14497\
        );

    \I__2111\ : InMux
    port map (
            O => \N__14502\,
            I => \N__14494\
        );

    \I__2110\ : InMux
    port map (
            O => \N__14501\,
            I => \N__14491\
        );

    \I__2109\ : InMux
    port map (
            O => \N__14500\,
            I => \N__14488\
        );

    \I__2108\ : Sp12to4
    port map (
            O => \N__14497\,
            I => \N__14483\
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__14494\,
            I => \N__14483\
        );

    \I__2106\ : LocalMux
    port map (
            O => \N__14491\,
            I => \N__14480\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__14488\,
            I => \N__14477\
        );

    \I__2104\ : Span12Mux_s5_v
    port map (
            O => \N__14483\,
            I => \N__14474\
        );

    \I__2103\ : Odrv4
    port map (
            O => \N__14480\,
            I => \Lab_UT.dictrl.currState_fast_0\
        );

    \I__2102\ : Odrv4
    port map (
            O => \N__14477\,
            I => \Lab_UT.dictrl.currState_fast_0\
        );

    \I__2101\ : Odrv12
    port map (
            O => \N__14474\,
            I => \Lab_UT.dictrl.currState_fast_0\
        );

    \I__2100\ : CascadeMux
    port map (
            O => \N__14467\,
            I => \Lab_UT.dictrl.g1_4_1_0_cascade_\
        );

    \I__2099\ : InMux
    port map (
            O => \N__14464\,
            I => \N__14461\
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__14461\,
            I => \Lab_UT.dictrl.de_littleA_0\
        );

    \I__2097\ : CascadeMux
    port map (
            O => \N__14458\,
            I => \Lab_UT.dictrl.g1_4_cascade_\
        );

    \I__2096\ : InMux
    port map (
            O => \N__14455\,
            I => \N__14452\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__14452\,
            I => \N__14449\
        );

    \I__2094\ : Span4Mux_v
    port map (
            O => \N__14449\,
            I => \N__14446\
        );

    \I__2093\ : Odrv4
    port map (
            O => \N__14446\,
            I => \Lab_UT.dictrl.N_17_0_0\
        );

    \I__2092\ : InMux
    port map (
            O => \N__14443\,
            I => \N__14440\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__14440\,
            I => \Lab_UT.dictrl.decoder.g0_5_1\
        );

    \I__2090\ : CascadeMux
    port map (
            O => \N__14437\,
            I => \N__14434\
        );

    \I__2089\ : InMux
    port map (
            O => \N__14434\,
            I => \N__14431\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__14431\,
            I => \Lab_UT.dictrl.m7_sx\
        );

    \I__2087\ : InMux
    port map (
            O => \N__14428\,
            I => \N__14424\
        );

    \I__2086\ : InMux
    port map (
            O => \N__14427\,
            I => \N__14421\
        );

    \I__2085\ : LocalMux
    port map (
            O => \N__14424\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_3\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__14421\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_3\
        );

    \I__2083\ : InMux
    port map (
            O => \N__14416\,
            I => \N__14410\
        );

    \I__2082\ : InMux
    port map (
            O => \N__14415\,
            I => \N__14407\
        );

    \I__2081\ : InMux
    port map (
            O => \N__14414\,
            I => \N__14402\
        );

    \I__2080\ : InMux
    port map (
            O => \N__14413\,
            I => \N__14402\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__14410\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_0\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__14407\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_0\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__14402\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_0\
        );

    \I__2076\ : InMux
    port map (
            O => \N__14395\,
            I => \N__14392\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__14392\,
            I => \buart.Z_rx.Z_baudgen.ser_clk_3\
        );

    \I__2074\ : InMux
    port map (
            O => \N__14389\,
            I => \N__14386\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__14386\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO\
        );

    \I__2072\ : CascadeMux
    port map (
            O => \N__14383\,
            I => \buart.Z_rx.ser_clk_cascade_\
        );

    \I__2071\ : CascadeMux
    port map (
            O => \N__14380\,
            I => \N__14376\
        );

    \I__2070\ : InMux
    port map (
            O => \N__14379\,
            I => \N__14372\
        );

    \I__2069\ : InMux
    port map (
            O => \N__14376\,
            I => \N__14367\
        );

    \I__2068\ : InMux
    port map (
            O => \N__14375\,
            I => \N__14367\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__14372\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_4\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__14367\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_4\
        );

    \I__2065\ : CascadeMux
    port map (
            O => \N__14362\,
            I => \N__14358\
        );

    \I__2064\ : InMux
    port map (
            O => \N__14361\,
            I => \N__14353\
        );

    \I__2063\ : InMux
    port map (
            O => \N__14358\,
            I => \N__14353\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__14353\,
            I => bu_rx_data_fast_7
        );

    \I__2061\ : CascadeMux
    port map (
            O => \N__14350\,
            I => \Lab_UT.dictrl.decoder.g0_5_0_cascade_\
        );

    \I__2060\ : InMux
    port map (
            O => \N__14347\,
            I => \N__14344\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__14344\,
            I => \N__14341\
        );

    \I__2058\ : Odrv4
    port map (
            O => \N__14341\,
            I => \Lab_UT.dictrl.de_cr_0_0\
        );

    \I__2057\ : InMux
    port map (
            O => \N__14338\,
            I => \N__14335\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__14335\,
            I => \N__14332\
        );

    \I__2055\ : Odrv4
    port map (
            O => \N__14332\,
            I => \Lab_UT.dictrl.decoder.g0_6_0\
        );

    \I__2054\ : InMux
    port map (
            O => \N__14329\,
            I => \N__14323\
        );

    \I__2053\ : InMux
    port map (
            O => \N__14328\,
            I => \N__14323\
        );

    \I__2052\ : LocalMux
    port map (
            O => \N__14323\,
            I => bu_rx_data_fast_6
        );

    \I__2051\ : InMux
    port map (
            O => \N__14320\,
            I => \N__14317\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__14317\,
            I => \Lab_UT.dictrl.decoder.g0Z0Z_4\
        );

    \I__2049\ : InMux
    port map (
            O => \N__14314\,
            I => \N__14308\
        );

    \I__2048\ : InMux
    port map (
            O => \N__14313\,
            I => \N__14308\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__14308\,
            I => bu_rx_data_fast_4
        );

    \I__2046\ : InMux
    port map (
            O => \N__14305\,
            I => \N__14299\
        );

    \I__2045\ : InMux
    port map (
            O => \N__14304\,
            I => \N__14299\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__14299\,
            I => bu_rx_data_fast_5
        );

    \I__2043\ : CascadeMux
    port map (
            O => \N__14296\,
            I => \N__14293\
        );

    \I__2042\ : InMux
    port map (
            O => \N__14293\,
            I => \N__14289\
        );

    \I__2041\ : InMux
    port map (
            O => \N__14292\,
            I => \N__14286\
        );

    \I__2040\ : LocalMux
    port map (
            O => \N__14289\,
            I => \N__14283\
        );

    \I__2039\ : LocalMux
    port map (
            O => \N__14286\,
            I => \N__14278\
        );

    \I__2038\ : Span4Mux_h
    port map (
            O => \N__14283\,
            I => \N__14278\
        );

    \I__2037\ : Odrv4
    port map (
            O => \N__14278\,
            I => \buart.Z_rx.hhZ0Z_0\
        );

    \I__2036\ : CascadeMux
    port map (
            O => \N__14275\,
            I => \buart.Z_rx.bitcount_fast_es_RNIAJ1GZ0Z_3_cascade_\
        );

    \I__2035\ : CascadeMux
    port map (
            O => \N__14272\,
            I => \bu_rx_data_rdy_cascade_\
        );

    \I__2034\ : CascadeMux
    port map (
            O => \N__14269\,
            I => \N__14265\
        );

    \I__2033\ : InMux
    port map (
            O => \N__14268\,
            I => \N__14262\
        );

    \I__2032\ : InMux
    port map (
            O => \N__14265\,
            I => \N__14259\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__14262\,
            I => \N__14256\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__14259\,
            I => \N__14253\
        );

    \I__2029\ : Span4Mux_h
    port map (
            O => \N__14256\,
            I => \N__14250\
        );

    \I__2028\ : Span4Mux_h
    port map (
            O => \N__14253\,
            I => \N__14247\
        );

    \I__2027\ : Odrv4
    port map (
            O => \N__14250\,
            I => \Lab_UT.dictrl.N_5_0_1\
        );

    \I__2026\ : Odrv4
    port map (
            O => \N__14247\,
            I => \Lab_UT.dictrl.N_5_0_1\
        );

    \I__2025\ : CascadeMux
    port map (
            O => \N__14242\,
            I => \Lab_UT.dictrl.g0_3_1_cascade_\
        );

    \I__2024\ : InMux
    port map (
            O => \N__14239\,
            I => \N__14236\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__14236\,
            I => \N__14233\
        );

    \I__2022\ : Odrv4
    port map (
            O => \N__14233\,
            I => \Lab_UT.dictrl.g0_1_0_0\
        );

    \I__2021\ : InMux
    port map (
            O => \N__14230\,
            I => \N__14227\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__14227\,
            I => bu_rx_data_fast_0
        );

    \I__2019\ : InMux
    port map (
            O => \N__14224\,
            I => \N__14219\
        );

    \I__2018\ : InMux
    port map (
            O => \N__14223\,
            I => \N__14214\
        );

    \I__2017\ : InMux
    port map (
            O => \N__14222\,
            I => \N__14214\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__14219\,
            I => \Lab_UT.dictrl.de_num_1_2\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__14214\,
            I => \Lab_UT.dictrl.de_num_1_2\
        );

    \I__2014\ : InMux
    port map (
            O => \N__14209\,
            I => \N__14206\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__14206\,
            I => \N__14202\
        );

    \I__2012\ : InMux
    port map (
            O => \N__14205\,
            I => \N__14199\
        );

    \I__2011\ : Odrv4
    port map (
            O => \N__14202\,
            I => \Lab_UT.dictrl.N_23_0_0\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__14199\,
            I => \Lab_UT.dictrl.N_23_0_0\
        );

    \I__2009\ : InMux
    port map (
            O => \N__14194\,
            I => \N__14191\
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__14191\,
            I => \Lab_UT.dictrl.N_13_0_0\
        );

    \I__2007\ : CascadeMux
    port map (
            O => \N__14188\,
            I => \Lab_UT.dictrl.N_14_0_0_0_cascade_\
        );

    \I__2006\ : InMux
    port map (
            O => \N__14185\,
            I => \N__14182\
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__14182\,
            I => \Lab_UT.dictrl.N_1609_0_0\
        );

    \I__2004\ : InMux
    port map (
            O => \N__14179\,
            I => \N__14176\
        );

    \I__2003\ : LocalMux
    port map (
            O => \N__14176\,
            I => \N__14172\
        );

    \I__2002\ : InMux
    port map (
            O => \N__14175\,
            I => \N__14169\
        );

    \I__2001\ : Span4Mux_v
    port map (
            O => \N__14172\,
            I => \N__14164\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__14169\,
            I => \N__14164\
        );

    \I__1999\ : Odrv4
    port map (
            O => \N__14164\,
            I => \Lab_UT.dictrl.N_8\
        );

    \I__1998\ : InMux
    port map (
            O => \N__14161\,
            I => \N__14157\
        );

    \I__1997\ : InMux
    port map (
            O => \N__14160\,
            I => \N__14153\
        );

    \I__1996\ : LocalMux
    port map (
            O => \N__14157\,
            I => \N__14150\
        );

    \I__1995\ : InMux
    port map (
            O => \N__14156\,
            I => \N__14147\
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__14153\,
            I => \Lab_UT.dictrl.N_7\
        );

    \I__1993\ : Odrv4
    port map (
            O => \N__14150\,
            I => \Lab_UT.dictrl.N_7\
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__14147\,
            I => \Lab_UT.dictrl.N_7\
        );

    \I__1991\ : CascadeMux
    port map (
            O => \N__14140\,
            I => \Lab_UT.dictrl.N_9_0_cascade_\
        );

    \I__1990\ : InMux
    port map (
            O => \N__14137\,
            I => \N__14134\
        );

    \I__1989\ : LocalMux
    port map (
            O => \N__14134\,
            I => \Lab_UT.dictrl.g0_6\
        );

    \I__1988\ : InMux
    port map (
            O => \N__14131\,
            I => \N__14128\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__14128\,
            I => \Lab_UT.dictrl.N_6_0\
        );

    \I__1986\ : InMux
    port map (
            O => \N__14125\,
            I => \N__14122\
        );

    \I__1985\ : LocalMux
    port map (
            O => \N__14122\,
            I => \N__14119\
        );

    \I__1984\ : Span4Mux_h
    port map (
            O => \N__14119\,
            I => \N__14116\
        );

    \I__1983\ : Odrv4
    port map (
            O => \N__14116\,
            I => \Lab_UT.dictrl.N_9\
        );

    \I__1982\ : InMux
    port map (
            O => \N__14113\,
            I => \N__14110\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__14110\,
            I => \Lab_UT.dictrl.m15_am\
        );

    \I__1980\ : InMux
    port map (
            O => \N__14107\,
            I => \N__14104\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__14104\,
            I => \Lab_UT.dictrl.N_20_1\
        );

    \I__1978\ : InMux
    port map (
            O => \N__14101\,
            I => \N__14098\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__14098\,
            I => \N__14092\
        );

    \I__1976\ : CascadeMux
    port map (
            O => \N__14097\,
            I => \N__14089\
        );

    \I__1975\ : CascadeMux
    port map (
            O => \N__14096\,
            I => \N__14084\
        );

    \I__1974\ : CascadeMux
    port map (
            O => \N__14095\,
            I => \N__14080\
        );

    \I__1973\ : Span4Mux_h
    port map (
            O => \N__14092\,
            I => \N__14077\
        );

    \I__1972\ : InMux
    port map (
            O => \N__14089\,
            I => \N__14064\
        );

    \I__1971\ : InMux
    port map (
            O => \N__14088\,
            I => \N__14064\
        );

    \I__1970\ : InMux
    port map (
            O => \N__14087\,
            I => \N__14064\
        );

    \I__1969\ : InMux
    port map (
            O => \N__14084\,
            I => \N__14064\
        );

    \I__1968\ : InMux
    port map (
            O => \N__14083\,
            I => \N__14064\
        );

    \I__1967\ : InMux
    port map (
            O => \N__14080\,
            I => \N__14064\
        );

    \I__1966\ : Odrv4
    port map (
            O => \N__14077\,
            I => \Lab_UT.dictrl.currState_0_rep1\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__14064\,
            I => \Lab_UT.dictrl.currState_0_rep1\
        );

    \I__1964\ : InMux
    port map (
            O => \N__14059\,
            I => \N__14056\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__14056\,
            I => \Lab_UT.dictrl.r_dicLdMtens17_1\
        );

    \I__1962\ : CascadeMux
    port map (
            O => \N__14053\,
            I => \N__14050\
        );

    \I__1961\ : InMux
    port map (
            O => \N__14050\,
            I => \N__14047\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__14047\,
            I => \N__14044\
        );

    \I__1959\ : Span4Mux_v
    port map (
            O => \N__14044\,
            I => \N__14041\
        );

    \I__1958\ : Odrv4
    port map (
            O => \N__14041\,
            I => \Lab_UT.dictrl.r_dicLdMtens22_2\
        );

    \I__1957\ : CascadeMux
    port map (
            O => \N__14038\,
            I => \Lab_UT.dictrl.N_34_cascade_\
        );

    \I__1956\ : InMux
    port map (
            O => \N__14035\,
            I => \N__14026\
        );

    \I__1955\ : InMux
    port map (
            O => \N__14034\,
            I => \N__14026\
        );

    \I__1954\ : InMux
    port map (
            O => \N__14033\,
            I => \N__14026\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__14026\,
            I => \N__14022\
        );

    \I__1952\ : InMux
    port map (
            O => \N__14025\,
            I => \N__14019\
        );

    \I__1951\ : Span4Mux_h
    port map (
            O => \N__14022\,
            I => \N__14016\
        );

    \I__1950\ : LocalMux
    port map (
            O => \N__14019\,
            I => \Lab_UT.dictrl.currState_2_RNI0P25DZ0Z_1\
        );

    \I__1949\ : Odrv4
    port map (
            O => \N__14016\,
            I => \Lab_UT.dictrl.currState_2_RNI0P25DZ0Z_1\
        );

    \I__1948\ : CascadeMux
    port map (
            O => \N__14011\,
            I => \Lab_UT.dictrl.m15_bm_cascade_\
        );

    \I__1947\ : CascadeMux
    port map (
            O => \N__14008\,
            I => \N__14004\
        );

    \I__1946\ : CascadeMux
    port map (
            O => \N__14007\,
            I => \N__14001\
        );

    \I__1945\ : InMux
    port map (
            O => \N__14004\,
            I => \N__13998\
        );

    \I__1944\ : InMux
    port map (
            O => \N__14001\,
            I => \N__13995\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__13998\,
            I => \N__13992\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__13995\,
            I => \Lab_UT.dictrl.nextState_0_0\
        );

    \I__1941\ : Odrv4
    port map (
            O => \N__13992\,
            I => \Lab_UT.dictrl.nextState_0_0\
        );

    \I__1940\ : InMux
    port map (
            O => \N__13987\,
            I => \N__13984\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__13984\,
            I => \Lab_UT.dictrl.N_7_0\
        );

    \I__1938\ : InMux
    port map (
            O => \N__13981\,
            I => \N__13978\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__13978\,
            I => \Lab_UT.dictrl.N_1609_1\
        );

    \I__1936\ : InMux
    port map (
            O => \N__13975\,
            I => \N__13971\
        );

    \I__1935\ : CascadeMux
    port map (
            O => \N__13974\,
            I => \N__13968\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__13971\,
            I => \N__13965\
        );

    \I__1933\ : InMux
    port map (
            O => \N__13968\,
            I => \N__13962\
        );

    \I__1932\ : Odrv4
    port map (
            O => \N__13965\,
            I => \Lab_UT.dictrl.N_38\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__13962\,
            I => \Lab_UT.dictrl.N_38\
        );

    \I__1930\ : InMux
    port map (
            O => \N__13957\,
            I => \N__13954\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__13954\,
            I => \Lab_UT.dictrl.currState_ret_5_RNOZ0Z_0\
        );

    \I__1928\ : CascadeMux
    port map (
            O => \N__13951\,
            I => \Lab_UT.dictrl.N_12_0_cascade_\
        );

    \I__1927\ : InMux
    port map (
            O => \N__13948\,
            I => \N__13945\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__13945\,
            I => \N__13942\
        );

    \I__1925\ : Odrv4
    port map (
            O => \N__13942\,
            I => \Lab_UT.dictrl.G_28_0_a5_2_1\
        );

    \I__1924\ : CascadeMux
    port map (
            O => \N__13939\,
            I => \N__13935\
        );

    \I__1923\ : InMux
    port map (
            O => \N__13938\,
            I => \N__13932\
        );

    \I__1922\ : InMux
    port map (
            O => \N__13935\,
            I => \N__13929\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__13932\,
            I => \N__13926\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__13929\,
            I => \Lab_UT.dictrl.dicLdAMtensZ0\
        );

    \I__1919\ : Odrv12
    port map (
            O => \N__13926\,
            I => \Lab_UT.dictrl.dicLdAMtensZ0\
        );

    \I__1918\ : InMux
    port map (
            O => \N__13921\,
            I => \N__13917\
        );

    \I__1917\ : InMux
    port map (
            O => \N__13920\,
            I => \N__13914\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__13917\,
            I => \Lab_UT.dictrl.dicLdAMtens_rst\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__13914\,
            I => \Lab_UT.dictrl.dicLdAMtens_rst\
        );

    \I__1914\ : InMux
    port map (
            O => \N__13909\,
            I => \N__13906\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__13906\,
            I => \Lab_UT.dictrl.r_dicLdMtens16_1\
        );

    \I__1912\ : CascadeMux
    port map (
            O => \N__13903\,
            I => \Lab_UT.dictrl.g0_10_0_N_4L6_1_cascade_\
        );

    \I__1911\ : SRMux
    port map (
            O => \N__13900\,
            I => \N__13897\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__13897\,
            I => \N__13893\
        );

    \I__1909\ : InMux
    port map (
            O => \N__13896\,
            I => \N__13890\
        );

    \I__1908\ : Span4Mux_h
    port map (
            O => \N__13893\,
            I => \N__13887\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__13890\,
            I => \N__13884\
        );

    \I__1906\ : Span4Mux_v
    port map (
            O => \N__13887\,
            I => \N__13881\
        );

    \I__1905\ : Span4Mux_h
    port map (
            O => \N__13884\,
            I => \N__13878\
        );

    \I__1904\ : Odrv4
    port map (
            O => \N__13881\,
            I => \Lab_UT.dictrl.currState_ret_RNI7FNUZ0\
        );

    \I__1903\ : Odrv4
    port map (
            O => \N__13878\,
            I => \Lab_UT.dictrl.currState_ret_RNI7FNUZ0\
        );

    \I__1902\ : CascadeMux
    port map (
            O => \N__13873\,
            I => \Lab_UT.Mone_at_0_cascade_\
        );

    \I__1901\ : InMux
    port map (
            O => \N__13870\,
            I => \N__13867\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__13867\,
            I => \Lab_UT.N_77_0\
        );

    \I__1899\ : InMux
    port map (
            O => \N__13864\,
            I => \N__13859\
        );

    \I__1898\ : InMux
    port map (
            O => \N__13863\,
            I => \N__13854\
        );

    \I__1897\ : InMux
    port map (
            O => \N__13862\,
            I => \N__13854\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__13859\,
            I => \N__13851\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__13854\,
            I => \N__13848\
        );

    \I__1894\ : Span4Mux_h
    port map (
            O => \N__13851\,
            I => \N__13845\
        );

    \I__1893\ : Span4Mux_h
    port map (
            O => \N__13848\,
            I => \N__13842\
        );

    \I__1892\ : Odrv4
    port map (
            O => \N__13845\,
            I => \Lab_UT.dictrl.N_23\
        );

    \I__1891\ : Odrv4
    port map (
            O => \N__13842\,
            I => \Lab_UT.dictrl.N_23\
        );

    \I__1890\ : CascadeMux
    port map (
            O => \N__13837\,
            I => \Lab_UT.dictrl.N_23_cascade_\
        );

    \I__1889\ : CascadeMux
    port map (
            O => \N__13834\,
            I => \N__13831\
        );

    \I__1888\ : InMux
    port map (
            O => \N__13831\,
            I => \N__13824\
        );

    \I__1887\ : InMux
    port map (
            O => \N__13830\,
            I => \N__13824\
        );

    \I__1886\ : InMux
    port map (
            O => \N__13829\,
            I => \N__13821\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__13824\,
            I => \N__13818\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__13821\,
            I => \N__13815\
        );

    \I__1883\ : Span4Mux_s3_h
    port map (
            O => \N__13818\,
            I => \N__13812\
        );

    \I__1882\ : Span4Mux_h
    port map (
            O => \N__13815\,
            I => \N__13809\
        );

    \I__1881\ : Odrv4
    port map (
            O => \N__13812\,
            I => \Lab_UT.dictrl.nextState_RNIA8EV3Z0Z_1\
        );

    \I__1880\ : Odrv4
    port map (
            O => \N__13809\,
            I => \Lab_UT.dictrl.nextState_RNIA8EV3Z0Z_1\
        );

    \I__1879\ : InMux
    port map (
            O => \N__13804\,
            I => \N__13801\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__13801\,
            I => \Lab_UT.dictrl.N_10\
        );

    \I__1877\ : CascadeMux
    port map (
            O => \N__13798\,
            I => \Lab_UT.segmentUQ_0_0_cascade_\
        );

    \I__1876\ : CascadeMux
    port map (
            O => \N__13795\,
            I => \Lab_UT.N_65_0_cascade_\
        );

    \I__1875\ : InMux
    port map (
            O => \N__13792\,
            I => \N__13789\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__13789\,
            I => \Lab_UT.segment_1_0_6\
        );

    \I__1873\ : CascadeMux
    port map (
            O => \N__13786\,
            I => \Lab_UT.N_76_0_cascade_\
        );

    \I__1872\ : InMux
    port map (
            O => \N__13783\,
            I => \N__13780\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__13780\,
            I => \uu2.bitmapZ0Z_72\
        );

    \I__1870\ : CascadeMux
    port map (
            O => \N__13777\,
            I => \N__13774\
        );

    \I__1869\ : InMux
    port map (
            O => \N__13774\,
            I => \N__13771\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__13771\,
            I => \uu2.bitmapZ0Z_200\
        );

    \I__1867\ : InMux
    port map (
            O => \N__13768\,
            I => \N__13765\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__13765\,
            I => \uu2.bitmap_RNIOS152Z0Z_72\
        );

    \I__1865\ : InMux
    port map (
            O => \N__13762\,
            I => \N__13759\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__13759\,
            I => \uu2.bitmapZ0Z_40\
        );

    \I__1863\ : CascadeMux
    port map (
            O => \N__13756\,
            I => \N__13753\
        );

    \I__1862\ : InMux
    port map (
            O => \N__13753\,
            I => \N__13750\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__13750\,
            I => \uu2.bitmapZ0Z_296\
        );

    \I__1860\ : CascadeMux
    port map (
            O => \N__13747\,
            I => \uu2.bitmap_pmux_25_am_1_cascade_\
        );

    \I__1859\ : InMux
    port map (
            O => \N__13744\,
            I => \N__13741\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__13741\,
            I => \N__13738\
        );

    \I__1857\ : Odrv4
    port map (
            O => \N__13738\,
            I => \uu2.bitmapZ0Z_197\
        );

    \I__1856\ : InMux
    port map (
            O => \N__13735\,
            I => \N__13732\
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__13732\,
            I => \uu2.bitmapZ0Z_66\
        );

    \I__1854\ : CascadeMux
    port map (
            O => \N__13729\,
            I => \uu2.bitmap_RNI2JA82Z0Z_212_cascade_\
        );

    \I__1853\ : InMux
    port map (
            O => \N__13726\,
            I => \N__13722\
        );

    \I__1852\ : InMux
    port map (
            O => \N__13725\,
            I => \N__13719\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__13722\,
            I => \uu2.N_31_i\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__13719\,
            I => \uu2.N_31_i\
        );

    \I__1849\ : InMux
    port map (
            O => \N__13714\,
            I => \N__13711\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__13711\,
            I => \uu2.bitmap_RNIM7D32Z0Z_69\
        );

    \I__1847\ : CascadeMux
    port map (
            O => \N__13708\,
            I => \uu2.bitmap_pmux_27_ns_1_cascade_\
        );

    \I__1846\ : InMux
    port map (
            O => \N__13705\,
            I => \N__13702\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__13702\,
            I => \uu2.N_407\
        );

    \I__1844\ : CascadeMux
    port map (
            O => \N__13699\,
            I => \uu2.un404_ci_0_cascade_\
        );

    \I__1843\ : CascadeMux
    port map (
            O => \N__13696\,
            I => \N__13693\
        );

    \I__1842\ : InMux
    port map (
            O => \N__13693\,
            I => \N__13689\
        );

    \I__1841\ : CascadeMux
    port map (
            O => \N__13692\,
            I => \N__13685\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__13689\,
            I => \N__13681\
        );

    \I__1839\ : InMux
    port map (
            O => \N__13688\,
            I => \N__13674\
        );

    \I__1838\ : InMux
    port map (
            O => \N__13685\,
            I => \N__13674\
        );

    \I__1837\ : InMux
    port map (
            O => \N__13684\,
            I => \N__13674\
        );

    \I__1836\ : Odrv4
    port map (
            O => \N__13681\,
            I => \uu2.r_addrZ0Z_6\
        );

    \I__1835\ : LocalMux
    port map (
            O => \N__13674\,
            I => \uu2.r_addrZ0Z_6\
        );

    \I__1834\ : CascadeMux
    port map (
            O => \N__13669\,
            I => \N__13666\
        );

    \I__1833\ : InMux
    port map (
            O => \N__13666\,
            I => \N__13663\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__13663\,
            I => \N__13659\
        );

    \I__1831\ : CascadeMux
    port map (
            O => \N__13662\,
            I => \N__13656\
        );

    \I__1830\ : Span4Mux_h
    port map (
            O => \N__13659\,
            I => \N__13651\
        );

    \I__1829\ : InMux
    port map (
            O => \N__13656\,
            I => \N__13648\
        );

    \I__1828\ : InMux
    port map (
            O => \N__13655\,
            I => \N__13643\
        );

    \I__1827\ : InMux
    port map (
            O => \N__13654\,
            I => \N__13643\
        );

    \I__1826\ : Odrv4
    port map (
            O => \N__13651\,
            I => \uu2.r_addrZ0Z_2\
        );

    \I__1825\ : LocalMux
    port map (
            O => \N__13648\,
            I => \uu2.r_addrZ0Z_2\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__13643\,
            I => \uu2.r_addrZ0Z_2\
        );

    \I__1823\ : CascadeMux
    port map (
            O => \N__13636\,
            I => \N__13633\
        );

    \I__1822\ : InMux
    port map (
            O => \N__13633\,
            I => \N__13630\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__13630\,
            I => \N__13627\
        );

    \I__1820\ : Span4Mux_h
    port map (
            O => \N__13627\,
            I => \N__13620\
        );

    \I__1819\ : InMux
    port map (
            O => \N__13626\,
            I => \N__13615\
        );

    \I__1818\ : InMux
    port map (
            O => \N__13625\,
            I => \N__13615\
        );

    \I__1817\ : InMux
    port map (
            O => \N__13624\,
            I => \N__13610\
        );

    \I__1816\ : InMux
    port map (
            O => \N__13623\,
            I => \N__13610\
        );

    \I__1815\ : Odrv4
    port map (
            O => \N__13620\,
            I => \uu2.r_addrZ0Z_1\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__13615\,
            I => \uu2.r_addrZ0Z_1\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__13610\,
            I => \uu2.r_addrZ0Z_1\
        );

    \I__1812\ : CascadeMux
    port map (
            O => \N__13603\,
            I => \N__13600\
        );

    \I__1811\ : InMux
    port map (
            O => \N__13600\,
            I => \N__13597\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__13597\,
            I => \N__13594\
        );

    \I__1809\ : Span4Mux_v
    port map (
            O => \N__13594\,
            I => \N__13590\
        );

    \I__1808\ : CascadeMux
    port map (
            O => \N__13593\,
            I => \N__13586\
        );

    \I__1807\ : Sp12to4
    port map (
            O => \N__13590\,
            I => \N__13580\
        );

    \I__1806\ : InMux
    port map (
            O => \N__13589\,
            I => \N__13573\
        );

    \I__1805\ : InMux
    port map (
            O => \N__13586\,
            I => \N__13573\
        );

    \I__1804\ : InMux
    port map (
            O => \N__13585\,
            I => \N__13573\
        );

    \I__1803\ : InMux
    port map (
            O => \N__13584\,
            I => \N__13568\
        );

    \I__1802\ : InMux
    port map (
            O => \N__13583\,
            I => \N__13568\
        );

    \I__1801\ : Odrv12
    port map (
            O => \N__13580\,
            I => \uu2.r_addrZ0Z_0\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__13573\,
            I => \uu2.r_addrZ0Z_0\
        );

    \I__1799\ : LocalMux
    port map (
            O => \N__13568\,
            I => \uu2.r_addrZ0Z_0\
        );

    \I__1798\ : CascadeMux
    port map (
            O => \N__13561\,
            I => \N__13558\
        );

    \I__1797\ : InMux
    port map (
            O => \N__13558\,
            I => \N__13553\
        );

    \I__1796\ : CascadeMux
    port map (
            O => \N__13557\,
            I => \N__13550\
        );

    \I__1795\ : CascadeMux
    port map (
            O => \N__13556\,
            I => \N__13547\
        );

    \I__1794\ : LocalMux
    port map (
            O => \N__13553\,
            I => \N__13544\
        );

    \I__1793\ : InMux
    port map (
            O => \N__13550\,
            I => \N__13539\
        );

    \I__1792\ : InMux
    port map (
            O => \N__13547\,
            I => \N__13539\
        );

    \I__1791\ : Odrv4
    port map (
            O => \N__13544\,
            I => \uu2.r_addrZ0Z_3\
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__13539\,
            I => \uu2.r_addrZ0Z_3\
        );

    \I__1789\ : CEMux
    port map (
            O => \N__13534\,
            I => \N__13531\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__13531\,
            I => \N__13528\
        );

    \I__1787\ : Odrv12
    port map (
            O => \N__13528\,
            I => \uu2.trig_rd_is_det_0\
        );

    \I__1786\ : CascadeMux
    port map (
            O => \N__13525\,
            I => \N__13522\
        );

    \I__1785\ : InMux
    port map (
            O => \N__13522\,
            I => \N__13519\
        );

    \I__1784\ : LocalMux
    port map (
            O => \N__13519\,
            I => \uu2.bitmap_pmux_sn_N_42\
        );

    \I__1783\ : CascadeMux
    port map (
            O => \N__13516\,
            I => \uu2.bitmap_pmux_26_bm_1_cascade_\
        );

    \I__1782\ : CascadeMux
    port map (
            O => \N__13513\,
            I => \N__13510\
        );

    \I__1781\ : InMux
    port map (
            O => \N__13510\,
            I => \N__13507\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__13507\,
            I => \uu2.N_161\
        );

    \I__1779\ : CascadeMux
    port map (
            O => \N__13504\,
            I => \uu2.N_400_cascade_\
        );

    \I__1778\ : InMux
    port map (
            O => \N__13501\,
            I => \N__13498\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__13498\,
            I => \uu2.N_409\
        );

    \I__1776\ : InMux
    port map (
            O => \N__13495\,
            I => \N__13492\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__13492\,
            I => \uu2.bitmap_RNI1PH82Z0Z_34\
        );

    \I__1774\ : InMux
    port map (
            O => \N__13489\,
            I => \N__13486\
        );

    \I__1773\ : LocalMux
    port map (
            O => \N__13486\,
            I => \uu2.N_404\
        );

    \I__1772\ : InMux
    port map (
            O => \N__13483\,
            I => \N__13480\
        );

    \I__1771\ : LocalMux
    port map (
            O => \N__13480\,
            I => \uu2.bitmapZ0Z_290\
        );

    \I__1770\ : CascadeMux
    port map (
            O => \N__13477\,
            I => \uu2.trig_rd_is_det_cascade_\
        );

    \I__1769\ : InMux
    port map (
            O => \N__13474\,
            I => \N__13471\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__13471\,
            I => \uu2.trig_rd_detZ0Z_1\
        );

    \I__1767\ : InMux
    port map (
            O => \N__13468\,
            I => \N__13463\
        );

    \I__1766\ : InMux
    port map (
            O => \N__13467\,
            I => \N__13460\
        );

    \I__1765\ : InMux
    port map (
            O => \N__13466\,
            I => \N__13457\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__13463\,
            I => \N__13454\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__13460\,
            I => \N__13451\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__13457\,
            I => \N__13447\
        );

    \I__1761\ : Span4Mux_v
    port map (
            O => \N__13454\,
            I => \N__13444\
        );

    \I__1760\ : Span4Mux_s2_v
    port map (
            O => \N__13451\,
            I => \N__13441\
        );

    \I__1759\ : InMux
    port map (
            O => \N__13450\,
            I => \N__13438\
        );

    \I__1758\ : Span4Mux_s3_h
    port map (
            O => \N__13447\,
            I => \N__13435\
        );

    \I__1757\ : Odrv4
    port map (
            O => \N__13444\,
            I => \uu2.vram_rd_clkZ0\
        );

    \I__1756\ : Odrv4
    port map (
            O => \N__13441\,
            I => \uu2.vram_rd_clkZ0\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__13438\,
            I => \uu2.vram_rd_clkZ0\
        );

    \I__1754\ : Odrv4
    port map (
            O => \N__13435\,
            I => \uu2.vram_rd_clkZ0\
        );

    \I__1753\ : InMux
    port map (
            O => \N__13426\,
            I => \N__13422\
        );

    \I__1752\ : InMux
    port map (
            O => \N__13425\,
            I => \N__13419\
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__13422\,
            I => \N__13416\
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__13419\,
            I => \N__13411\
        );

    \I__1749\ : Span4Mux_h
    port map (
            O => \N__13416\,
            I => \N__13411\
        );

    \I__1748\ : Odrv4
    port map (
            O => \N__13411\,
            I => \uu2.un1_l_count_1_0\
        );

    \I__1747\ : InMux
    port map (
            O => \N__13408\,
            I => \N__13402\
        );

    \I__1746\ : InMux
    port map (
            O => \N__13407\,
            I => \N__13402\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__13402\,
            I => \uu2.trig_rd_detZ0Z_0\
        );

    \I__1744\ : InMux
    port map (
            O => \N__13399\,
            I => \N__13396\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__13396\,
            I => \uu2.vbuf_raddr.un448_ci_0\
        );

    \I__1742\ : CascadeMux
    port map (
            O => \N__13393\,
            I => \uu2.vbuf_raddr.un426_ci_3_cascade_\
        );

    \I__1741\ : CascadeMux
    port map (
            O => \N__13390\,
            I => \N__13387\
        );

    \I__1740\ : InMux
    port map (
            O => \N__13387\,
            I => \N__13384\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__13384\,
            I => \N__13380\
        );

    \I__1738\ : InMux
    port map (
            O => \N__13383\,
            I => \N__13377\
        );

    \I__1737\ : Span4Mux_s3_h
    port map (
            O => \N__13380\,
            I => \N__13372\
        );

    \I__1736\ : LocalMux
    port map (
            O => \N__13377\,
            I => \N__13372\
        );

    \I__1735\ : Odrv4
    port map (
            O => \N__13372\,
            I => \uu2.r_addrZ0Z_8\
        );

    \I__1734\ : InMux
    port map (
            O => \N__13369\,
            I => \N__13366\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__13366\,
            I => \uu2.vbuf_raddr.un426_ci_3\
        );

    \I__1732\ : CascadeMux
    port map (
            O => \N__13363\,
            I => \N__13360\
        );

    \I__1731\ : InMux
    port map (
            O => \N__13360\,
            I => \N__13357\
        );

    \I__1730\ : LocalMux
    port map (
            O => \N__13357\,
            I => \N__13352\
        );

    \I__1729\ : InMux
    port map (
            O => \N__13356\,
            I => \N__13349\
        );

    \I__1728\ : InMux
    port map (
            O => \N__13355\,
            I => \N__13346\
        );

    \I__1727\ : Odrv4
    port map (
            O => \N__13352\,
            I => \uu2.r_addrZ0Z_7\
        );

    \I__1726\ : LocalMux
    port map (
            O => \N__13349\,
            I => \uu2.r_addrZ0Z_7\
        );

    \I__1725\ : LocalMux
    port map (
            O => \N__13346\,
            I => \uu2.r_addrZ0Z_7\
        );

    \I__1724\ : InMux
    port map (
            O => \N__13339\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_2\
        );

    \I__1723\ : InMux
    port map (
            O => \N__13336\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_3\
        );

    \I__1722\ : InMux
    port map (
            O => \N__13333\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_4\
        );

    \I__1721\ : CascadeMux
    port map (
            O => \N__13330\,
            I => \N__13326\
        );

    \I__1720\ : InMux
    port map (
            O => \N__13329\,
            I => \N__13321\
        );

    \I__1719\ : InMux
    port map (
            O => \N__13326\,
            I => \N__13321\
        );

    \I__1718\ : LocalMux
    port map (
            O => \N__13321\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_5\
        );

    \I__1717\ : CascadeMux
    port map (
            O => \N__13318\,
            I => \N__13315\
        );

    \I__1716\ : InMux
    port map (
            O => \N__13315\,
            I => \N__13312\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__13312\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO\
        );

    \I__1714\ : InMux
    port map (
            O => \N__13309\,
            I => \N__13300\
        );

    \I__1713\ : InMux
    port map (
            O => \N__13308\,
            I => \N__13300\
        );

    \I__1712\ : InMux
    port map (
            O => \N__13307\,
            I => \N__13300\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__13300\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_2\
        );

    \I__1710\ : CascadeMux
    port map (
            O => \N__13297\,
            I => \N__13293\
        );

    \I__1709\ : InMux
    port map (
            O => \N__13296\,
            I => \N__13285\
        );

    \I__1708\ : InMux
    port map (
            O => \N__13293\,
            I => \N__13285\
        );

    \I__1707\ : InMux
    port map (
            O => \N__13292\,
            I => \N__13285\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__13285\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_1\
        );

    \I__1705\ : CascadeMux
    port map (
            O => \N__13282\,
            I => \G_28_0_a5_0_4_cascade_\
        );

    \I__1704\ : CascadeMux
    port map (
            O => \N__13279\,
            I => \N__13276\
        );

    \I__1703\ : InMux
    port map (
            O => \N__13276\,
            I => \N__13273\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__13273\,
            I => \N__13270\
        );

    \I__1701\ : Odrv12
    port map (
            O => \N__13270\,
            I => \shifter_RNI1D8L1_4\
        );

    \I__1700\ : InMux
    port map (
            O => \N__13267\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_1\
        );

    \I__1699\ : CascadeMux
    port map (
            O => \N__13264\,
            I => \Lab_UT.dictrl.decoder.g0Z0Z_5_cascade_\
        );

    \I__1698\ : InMux
    port map (
            O => \N__13261\,
            I => \N__13258\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__13258\,
            I => \Lab_UT.dictrl.decoder.g0Z0Z_1\
        );

    \I__1696\ : CascadeMux
    port map (
            O => \N__13255\,
            I => \Lab_UT.dictrl.N_36_1_cascade_\
        );

    \I__1695\ : InMux
    port map (
            O => \N__13252\,
            I => \N__13249\
        );

    \I__1694\ : LocalMux
    port map (
            O => \N__13249\,
            I => \N__13246\
        );

    \I__1693\ : Odrv4
    port map (
            O => \N__13246\,
            I => \Lab_UT.dictrl.g1_0_1\
        );

    \I__1692\ : InMux
    port map (
            O => \N__13243\,
            I => \N__13240\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__13240\,
            I => \Lab_UT.dictrl.N_7_1\
        );

    \I__1690\ : CascadeMux
    port map (
            O => \N__13237\,
            I => \N__13234\
        );

    \I__1689\ : InMux
    port map (
            O => \N__13234\,
            I => \N__13230\
        );

    \I__1688\ : InMux
    port map (
            O => \N__13233\,
            I => \N__13227\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__13230\,
            I => \N__13224\
        );

    \I__1686\ : LocalMux
    port map (
            O => \N__13227\,
            I => \N__13220\
        );

    \I__1685\ : Span4Mux_h
    port map (
            O => \N__13224\,
            I => \N__13217\
        );

    \I__1684\ : InMux
    port map (
            O => \N__13223\,
            I => \N__13213\
        );

    \I__1683\ : Span4Mux_h
    port map (
            O => \N__13220\,
            I => \N__13210\
        );

    \I__1682\ : Span4Mux_s0_h
    port map (
            O => \N__13217\,
            I => \N__13207\
        );

    \I__1681\ : InMux
    port map (
            O => \N__13216\,
            I => \N__13204\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__13213\,
            I => \Lab_UT.dictrl.nextState_0_1\
        );

    \I__1679\ : Odrv4
    port map (
            O => \N__13210\,
            I => \Lab_UT.dictrl.nextState_0_1\
        );

    \I__1678\ : Odrv4
    port map (
            O => \N__13207\,
            I => \Lab_UT.dictrl.nextState_0_1\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__13204\,
            I => \Lab_UT.dictrl.nextState_0_1\
        );

    \I__1676\ : CascadeMux
    port map (
            O => \N__13195\,
            I => \Lab_UT.dictrl.N_20_cascade_\
        );

    \I__1675\ : InMux
    port map (
            O => \N__13192\,
            I => \N__13186\
        );

    \I__1674\ : InMux
    port map (
            O => \N__13191\,
            I => \N__13186\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__13186\,
            I => \Lab_UT.dictrl.G_28_0_a5_1\
        );

    \I__1672\ : InMux
    port map (
            O => \N__13183\,
            I => \N__13177\
        );

    \I__1671\ : InMux
    port map (
            O => \N__13182\,
            I => \N__13177\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__13177\,
            I => \Lab_UT.dictrl.N_19_0\
        );

    \I__1669\ : CascadeMux
    port map (
            O => \N__13174\,
            I => \Lab_UT.dictrl.N_8_3_cascade_\
        );

    \I__1668\ : CascadeMux
    port map (
            O => \N__13171\,
            I => \Lab_UT.dictrl.currState_2_0_rep2_RNIBGCIZ0Z9_cascade_\
        );

    \I__1667\ : InMux
    port map (
            O => \N__13168\,
            I => \N__13162\
        );

    \I__1666\ : InMux
    port map (
            O => \N__13167\,
            I => \N__13162\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__13162\,
            I => \Lab_UT.dictrl.G_28_0_0\
        );

    \I__1664\ : InMux
    port map (
            O => \N__13159\,
            I => \N__13156\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__13156\,
            I => \Lab_UT.dictrl.currState_2_0_rep2_RNIKH8PZ0Z2\
        );

    \I__1662\ : InMux
    port map (
            O => \N__13153\,
            I => \N__13150\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__13150\,
            I => \shifter_RNIS6CF1_5\
        );

    \I__1660\ : CascadeMux
    port map (
            O => \N__13147\,
            I => \Lab_UT.dictrl.m21_rn_1_0_cascade_\
        );

    \I__1659\ : InMux
    port map (
            O => \N__13144\,
            I => \N__13141\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__13141\,
            I => \Lab_UT.dictrl.m21_rn_0\
        );

    \I__1657\ : CascadeMux
    port map (
            O => \N__13138\,
            I => \Lab_UT.dictrl.g0_0_0_cascade_\
        );

    \I__1656\ : CascadeMux
    port map (
            O => \N__13135\,
            I => \Lab_UT.dictrl.N_1611_0_cascade_\
        );

    \I__1655\ : InMux
    port map (
            O => \N__13132\,
            I => \N__13129\
        );

    \I__1654\ : LocalMux
    port map (
            O => \N__13129\,
            I => \Lab_UT.dictrl.N_23_0\
        );

    \I__1653\ : CascadeMux
    port map (
            O => \N__13126\,
            I => \N__13123\
        );

    \I__1652\ : InMux
    port map (
            O => \N__13123\,
            I => \N__13120\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__13120\,
            I => \Lab_UT.dictrl.N_8_3\
        );

    \I__1650\ : InMux
    port map (
            O => \N__13117\,
            I => \N__13106\
        );

    \I__1649\ : InMux
    port map (
            O => \N__13116\,
            I => \N__13106\
        );

    \I__1648\ : InMux
    port map (
            O => \N__13115\,
            I => \N__13106\
        );

    \I__1647\ : InMux
    port map (
            O => \N__13114\,
            I => \N__13103\
        );

    \I__1646\ : InMux
    port map (
            O => \N__13113\,
            I => \N__13100\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__13106\,
            I => \N__13097\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__13103\,
            I => \uu2.l_countZ0Z_1\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__13100\,
            I => \uu2.l_countZ0Z_1\
        );

    \I__1642\ : Odrv4
    port map (
            O => \N__13097\,
            I => \uu2.l_countZ0Z_1\
        );

    \I__1641\ : CascadeMux
    port map (
            O => \N__13090\,
            I => \N__13085\
        );

    \I__1640\ : InMux
    port map (
            O => \N__13089\,
            I => \N__13080\
        );

    \I__1639\ : InMux
    port map (
            O => \N__13088\,
            I => \N__13080\
        );

    \I__1638\ : InMux
    port map (
            O => \N__13085\,
            I => \N__13074\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__13080\,
            I => \N__13071\
        );

    \I__1636\ : InMux
    port map (
            O => \N__13079\,
            I => \N__13066\
        );

    \I__1635\ : InMux
    port map (
            O => \N__13078\,
            I => \N__13066\
        );

    \I__1634\ : InMux
    port map (
            O => \N__13077\,
            I => \N__13063\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__13074\,
            I => \N__13060\
        );

    \I__1632\ : Span4Mux_h
    port map (
            O => \N__13071\,
            I => \N__13057\
        );

    \I__1631\ : LocalMux
    port map (
            O => \N__13066\,
            I => \uu2.l_countZ0Z_0\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__13063\,
            I => \uu2.l_countZ0Z_0\
        );

    \I__1629\ : Odrv4
    port map (
            O => \N__13060\,
            I => \uu2.l_countZ0Z_0\
        );

    \I__1628\ : Odrv4
    port map (
            O => \N__13057\,
            I => \uu2.l_countZ0Z_0\
        );

    \I__1627\ : CascadeMux
    port map (
            O => \N__13048\,
            I => \N__13045\
        );

    \I__1626\ : InMux
    port map (
            O => \N__13045\,
            I => \N__13039\
        );

    \I__1625\ : InMux
    port map (
            O => \N__13044\,
            I => \N__13039\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__13039\,
            I => \N__13036\
        );

    \I__1623\ : Span4Mux_s3_h
    port map (
            O => \N__13036\,
            I => \N__13033\
        );

    \I__1622\ : Odrv4
    port map (
            O => \N__13033\,
            I => \uu2.un284_ci\
        );

    \I__1621\ : CascadeMux
    port map (
            O => \N__13030\,
            I => \Lab_UT.dictrl.N_9_cascade_\
        );

    \I__1620\ : CascadeMux
    port map (
            O => \N__13027\,
            I => \Lab_UT.dictrl.N_21_1_cascade_\
        );

    \I__1619\ : InMux
    port map (
            O => \N__13024\,
            I => \N__13018\
        );

    \I__1618\ : InMux
    port map (
            O => \N__13023\,
            I => \N__13018\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__13018\,
            I => \N__13015\
        );

    \I__1616\ : Odrv4
    port map (
            O => \N__13015\,
            I => \uu2.w_data_displaying_2_i_a2_i_a3_1_0\
        );

    \I__1615\ : InMux
    port map (
            O => \N__13012\,
            I => \N__13008\
        );

    \I__1614\ : InMux
    port map (
            O => \N__13011\,
            I => \N__13004\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__13008\,
            I => \N__13001\
        );

    \I__1612\ : InMux
    port map (
            O => \N__13007\,
            I => \N__12998\
        );

    \I__1611\ : LocalMux
    port map (
            O => \N__13004\,
            I => \N__12995\
        );

    \I__1610\ : Span4Mux_v
    port map (
            O => \N__13001\,
            I => \N__12990\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__12998\,
            I => \N__12990\
        );

    \I__1608\ : Span4Mux_h
    port map (
            O => \N__12995\,
            I => \N__12978\
        );

    \I__1607\ : Span4Mux_v
    port map (
            O => \N__12990\,
            I => \N__12975\
        );

    \I__1606\ : InMux
    port map (
            O => \N__12989\,
            I => \N__12968\
        );

    \I__1605\ : InMux
    port map (
            O => \N__12988\,
            I => \N__12968\
        );

    \I__1604\ : InMux
    port map (
            O => \N__12987\,
            I => \N__12968\
        );

    \I__1603\ : InMux
    port map (
            O => \N__12986\,
            I => \N__12963\
        );

    \I__1602\ : InMux
    port map (
            O => \N__12985\,
            I => \N__12963\
        );

    \I__1601\ : InMux
    port map (
            O => \N__12984\,
            I => \N__12954\
        );

    \I__1600\ : InMux
    port map (
            O => \N__12983\,
            I => \N__12954\
        );

    \I__1599\ : InMux
    port map (
            O => \N__12982\,
            I => \N__12954\
        );

    \I__1598\ : InMux
    port map (
            O => \N__12981\,
            I => \N__12954\
        );

    \I__1597\ : Span4Mux_v
    port map (
            O => \N__12978\,
            I => \N__12951\
        );

    \I__1596\ : Odrv4
    port map (
            O => \N__12975\,
            I => \uu0.un4_l_count_0\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__12968\,
            I => \uu0.un4_l_count_0\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__12963\,
            I => \uu0.un4_l_count_0\
        );

    \I__1593\ : LocalMux
    port map (
            O => \N__12954\,
            I => \uu0.un4_l_count_0\
        );

    \I__1592\ : Odrv4
    port map (
            O => \N__12951\,
            I => \uu0.un4_l_count_0\
        );

    \I__1591\ : InMux
    port map (
            O => \N__12940\,
            I => \N__12935\
        );

    \I__1590\ : InMux
    port map (
            O => \N__12939\,
            I => \N__12932\
        );

    \I__1589\ : InMux
    port map (
            O => \N__12938\,
            I => \N__12929\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__12935\,
            I => \N__12926\
        );

    \I__1587\ : LocalMux
    port map (
            O => \N__12932\,
            I => \uu2.un1_l_count_2_0\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__12929\,
            I => \uu2.un1_l_count_2_0\
        );

    \I__1585\ : Odrv4
    port map (
            O => \N__12926\,
            I => \uu2.un1_l_count_2_0\
        );

    \I__1584\ : InMux
    port map (
            O => \N__12919\,
            I => \N__12916\
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__12916\,
            I => \N__12912\
        );

    \I__1582\ : InMux
    port map (
            O => \N__12915\,
            I => \N__12909\
        );

    \I__1581\ : Span4Mux_h
    port map (
            O => \N__12912\,
            I => \N__12906\
        );

    \I__1580\ : LocalMux
    port map (
            O => \N__12909\,
            I => \N__12903\
        );

    \I__1579\ : Span4Mux_v
    port map (
            O => \N__12906\,
            I => \N__12900\
        );

    \I__1578\ : Span4Mux_h
    port map (
            O => \N__12903\,
            I => \N__12897\
        );

    \I__1577\ : Odrv4
    port map (
            O => \N__12900\,
            I => \uu0.delay_lineZ0Z_0\
        );

    \I__1576\ : Odrv4
    port map (
            O => \N__12897\,
            I => \uu0.delay_lineZ0Z_0\
        );

    \I__1575\ : InMux
    port map (
            O => \N__12892\,
            I => \N__12889\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__12889\,
            I => \N__12886\
        );

    \I__1573\ : Odrv12
    port map (
            O => \N__12886\,
            I => \uu0.delay_lineZ0Z_1\
        );

    \I__1572\ : InMux
    port map (
            O => \N__12883\,
            I => \N__12880\
        );

    \I__1571\ : LocalMux
    port map (
            O => \N__12880\,
            I => \uu2.bitmap_pmux_sn_i7_mux_0\
        );

    \I__1570\ : CascadeMux
    port map (
            O => \N__12877\,
            I => \uu2.bitmap_pmux_29_0_cascade_\
        );

    \I__1569\ : CascadeMux
    port map (
            O => \N__12874\,
            I => \N__12871\
        );

    \I__1568\ : InMux
    port map (
            O => \N__12871\,
            I => \N__12865\
        );

    \I__1567\ : InMux
    port map (
            O => \N__12870\,
            I => \N__12865\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__12865\,
            I => \uu2.bitmap_pmux\
        );

    \I__1565\ : InMux
    port map (
            O => \N__12862\,
            I => \N__12859\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__12859\,
            I => \uu2.bitmap_pmux_sn_N_36\
        );

    \I__1563\ : InMux
    port map (
            O => \N__12856\,
            I => \N__12853\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__12853\,
            I => \N__12850\
        );

    \I__1561\ : Span4Mux_h
    port map (
            O => \N__12850\,
            I => \N__12847\
        );

    \I__1560\ : Odrv4
    port map (
            O => \N__12847\,
            I => vbuf_tx_data_6
        );

    \I__1559\ : InMux
    port map (
            O => \N__12844\,
            I => \N__12841\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__12841\,
            I => \N__12838\
        );

    \I__1557\ : Span4Mux_v
    port map (
            O => \N__12838\,
            I => \N__12835\
        );

    \I__1556\ : Odrv4
    port map (
            O => \N__12835\,
            I => \buart.Z_tx.shifterZ0Z_7\
        );

    \I__1555\ : CascadeMux
    port map (
            O => \N__12832\,
            I => \N__12827\
        );

    \I__1554\ : InMux
    port map (
            O => \N__12831\,
            I => \N__12820\
        );

    \I__1553\ : InMux
    port map (
            O => \N__12830\,
            I => \N__12820\
        );

    \I__1552\ : InMux
    port map (
            O => \N__12827\,
            I => \N__12808\
        );

    \I__1551\ : InMux
    port map (
            O => \N__12826\,
            I => \N__12803\
        );

    \I__1550\ : InMux
    port map (
            O => \N__12825\,
            I => \N__12803\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__12820\,
            I => \N__12800\
        );

    \I__1548\ : InMux
    port map (
            O => \N__12819\,
            I => \N__12781\
        );

    \I__1547\ : InMux
    port map (
            O => \N__12818\,
            I => \N__12781\
        );

    \I__1546\ : InMux
    port map (
            O => \N__12817\,
            I => \N__12781\
        );

    \I__1545\ : InMux
    port map (
            O => \N__12816\,
            I => \N__12781\
        );

    \I__1544\ : InMux
    port map (
            O => \N__12815\,
            I => \N__12781\
        );

    \I__1543\ : InMux
    port map (
            O => \N__12814\,
            I => \N__12781\
        );

    \I__1542\ : InMux
    port map (
            O => \N__12813\,
            I => \N__12781\
        );

    \I__1541\ : InMux
    port map (
            O => \N__12812\,
            I => \N__12781\
        );

    \I__1540\ : InMux
    port map (
            O => \N__12811\,
            I => \N__12778\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__12808\,
            I => \N__12771\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__12803\,
            I => \N__12771\
        );

    \I__1537\ : Span4Mux_h
    port map (
            O => \N__12800\,
            I => \N__12771\
        );

    \I__1536\ : InMux
    port map (
            O => \N__12799\,
            I => \N__12766\
        );

    \I__1535\ : InMux
    port map (
            O => \N__12798\,
            I => \N__12766\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__12781\,
            I => vbuf_tx_data_rdy
        );

    \I__1533\ : LocalMux
    port map (
            O => \N__12778\,
            I => vbuf_tx_data_rdy
        );

    \I__1532\ : Odrv4
    port map (
            O => \N__12771\,
            I => vbuf_tx_data_rdy
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__12766\,
            I => vbuf_tx_data_rdy
        );

    \I__1530\ : InMux
    port map (
            O => \N__12757\,
            I => \N__12754\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__12754\,
            I => \N__12751\
        );

    \I__1528\ : Span4Mux_v
    port map (
            O => \N__12751\,
            I => \N__12748\
        );

    \I__1527\ : Odrv4
    port map (
            O => \N__12748\,
            I => vbuf_tx_data_7
        );

    \I__1526\ : CascadeMux
    port map (
            O => \N__12745\,
            I => \N__12742\
        );

    \I__1525\ : InMux
    port map (
            O => \N__12742\,
            I => \N__12739\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__12739\,
            I => \buart.Z_tx.shifterZ0Z_8\
        );

    \I__1523\ : CEMux
    port map (
            O => \N__12736\,
            I => \N__12733\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__12733\,
            I => \N__12730\
        );

    \I__1521\ : Span4Mux_h
    port map (
            O => \N__12730\,
            I => \N__12726\
        );

    \I__1520\ : CEMux
    port map (
            O => \N__12729\,
            I => \N__12723\
        );

    \I__1519\ : Span4Mux_s0_h
    port map (
            O => \N__12726\,
            I => \N__12720\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__12723\,
            I => \N__12717\
        );

    \I__1517\ : Odrv4
    port map (
            O => \N__12720\,
            I => \buart.Z_tx.un1_uart_wr_i_0_i\
        );

    \I__1516\ : Odrv4
    port map (
            O => \N__12717\,
            I => \buart.Z_tx.un1_uart_wr_i_0_i\
        );

    \I__1515\ : IoInMux
    port map (
            O => \N__12712\,
            I => \N__12709\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__12709\,
            I => \N__12706\
        );

    \I__1513\ : Span4Mux_s3_h
    port map (
            O => \N__12706\,
            I => \N__12703\
        );

    \I__1512\ : Odrv4
    port map (
            O => \N__12703\,
            I => \uu0.un11_l_count_i\
        );

    \I__1511\ : CascadeMux
    port map (
            O => \N__12700\,
            I => \N__12697\
        );

    \I__1510\ : InMux
    port map (
            O => \N__12697\,
            I => \N__12694\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__12694\,
            I => \N__12691\
        );

    \I__1508\ : Span4Mux_s3_v
    port map (
            O => \N__12691\,
            I => \N__12688\
        );

    \I__1507\ : Odrv4
    port map (
            O => \N__12688\,
            I => \uu2.mem0.w_addr_7\
        );

    \I__1506\ : CascadeMux
    port map (
            O => \N__12685\,
            I => \N__12682\
        );

    \I__1505\ : InMux
    port map (
            O => \N__12682\,
            I => \N__12679\
        );

    \I__1504\ : LocalMux
    port map (
            O => \N__12679\,
            I => \N__12676\
        );

    \I__1503\ : Span4Mux_v
    port map (
            O => \N__12676\,
            I => \N__12673\
        );

    \I__1502\ : Odrv4
    port map (
            O => \N__12673\,
            I => \uu2.mem0.w_addr_1\
        );

    \I__1501\ : CascadeMux
    port map (
            O => \N__12670\,
            I => \uu2.N_51_cascade_\
        );

    \I__1500\ : InMux
    port map (
            O => \N__12667\,
            I => \N__12661\
        );

    \I__1499\ : InMux
    port map (
            O => \N__12666\,
            I => \N__12661\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__12661\,
            I => \uu2.N_34\
        );

    \I__1497\ : CascadeMux
    port map (
            O => \N__12658\,
            I => \uu2.N_34_cascade_\
        );

    \I__1496\ : InMux
    port map (
            O => \N__12655\,
            I => \N__12652\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__12652\,
            I => \uu2.mem0.w_data_0\
        );

    \I__1494\ : CascadeMux
    port map (
            O => \N__12649\,
            I => \uu2.bitmap_pmux_sn_m15_0_ns_1_cascade_\
        );

    \I__1493\ : InMux
    port map (
            O => \N__12646\,
            I => \N__12643\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__12643\,
            I => \uu2.bitmap_pmux_sn_N_65\
        );

    \I__1491\ : CascadeMux
    port map (
            O => \N__12640\,
            I => \uu2.bitmap_pmux_sn_m24_0_ns_1_cascade_\
        );

    \I__1490\ : CascadeMux
    port map (
            O => \N__12637\,
            I => \uu2.bitmap_pmux_sn_i5_mux_cascade_\
        );

    \I__1489\ : CascadeMux
    port map (
            O => \N__12634\,
            I => \N__12631\
        );

    \I__1488\ : InMux
    port map (
            O => \N__12631\,
            I => \N__12628\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__12628\,
            I => \uu2.mem0.w_addr_8\
        );

    \I__1486\ : InMux
    port map (
            O => \N__12625\,
            I => \N__12622\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__12622\,
            I => \N__12619\
        );

    \I__1484\ : Span4Mux_h
    port map (
            O => \N__12619\,
            I => \N__12616\
        );

    \I__1483\ : Odrv4
    port map (
            O => \N__12616\,
            I => \uu2.vram_rd_clk_detZ0Z_1\
        );

    \I__1482\ : InMux
    port map (
            O => \N__12613\,
            I => \N__12610\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__12610\,
            I => \N__12606\
        );

    \I__1480\ : InMux
    port map (
            O => \N__12609\,
            I => \N__12603\
        );

    \I__1479\ : Span4Mux_h
    port map (
            O => \N__12606\,
            I => \N__12600\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__12603\,
            I => \uu2.vram_rd_clk_detZ0Z_0\
        );

    \I__1477\ : Odrv4
    port map (
            O => \N__12600\,
            I => \uu2.vram_rd_clk_detZ0Z_0\
        );

    \I__1476\ : CEMux
    port map (
            O => \N__12595\,
            I => \N__12592\
        );

    \I__1475\ : LocalMux
    port map (
            O => \N__12592\,
            I => \N__12589\
        );

    \I__1474\ : Span4Mux_v
    port map (
            O => \N__12589\,
            I => \N__12586\
        );

    \I__1473\ : Span4Mux_s1_h
    port map (
            O => \N__12586\,
            I => \N__12583\
        );

    \I__1472\ : Odrv4
    port map (
            O => \N__12583\,
            I => \uu2.vram_rd_clk_det_RNI95711Z0Z_1\
        );

    \I__1471\ : InMux
    port map (
            O => \N__12580\,
            I => \N__12577\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__12577\,
            I => \uu2.mem0.w_data_4\
        );

    \I__1469\ : InMux
    port map (
            O => \N__12574\,
            I => \N__12571\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__12571\,
            I => \uu2.mem0.w_data_5\
        );

    \I__1467\ : InMux
    port map (
            O => \N__12568\,
            I => \N__12565\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__12565\,
            I => \uu2.N_37\
        );

    \I__1465\ : CascadeMux
    port map (
            O => \N__12562\,
            I => \uu2.N_37_cascade_\
        );

    \I__1464\ : InMux
    port map (
            O => \N__12559\,
            I => \N__12556\
        );

    \I__1463\ : LocalMux
    port map (
            O => \N__12556\,
            I => \uu2.mem0.w_data_3\
        );

    \I__1462\ : InMux
    port map (
            O => \N__12553\,
            I => \N__12550\
        );

    \I__1461\ : LocalMux
    port map (
            O => \N__12550\,
            I => \uu2.mem0.w_data_1\
        );

    \I__1460\ : InMux
    port map (
            O => \N__12547\,
            I => \N__12544\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__12544\,
            I => \Lab_UT.dictrl.G_19_0_a7_3_2\
        );

    \I__1458\ : InMux
    port map (
            O => \N__12541\,
            I => \N__12538\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__12538\,
            I => \G_19_0_a7_4_8\
        );

    \I__1456\ : InMux
    port map (
            O => \N__12535\,
            I => \N__12532\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__12532\,
            I => \G_19_0_a7_4_1\
        );

    \I__1454\ : CascadeMux
    port map (
            O => \N__12529\,
            I => \N__12526\
        );

    \I__1453\ : InMux
    port map (
            O => \N__12526\,
            I => \N__12514\
        );

    \I__1452\ : InMux
    port map (
            O => \N__12525\,
            I => \N__12514\
        );

    \I__1451\ : InMux
    port map (
            O => \N__12524\,
            I => \N__12514\
        );

    \I__1450\ : InMux
    port map (
            O => \N__12523\,
            I => \N__12514\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__12514\,
            I => \N__12509\
        );

    \I__1448\ : InMux
    port map (
            O => \N__12513\,
            I => \N__12506\
        );

    \I__1447\ : InMux
    port map (
            O => \N__12512\,
            I => \N__12503\
        );

    \I__1446\ : Span4Mux_v
    port map (
            O => \N__12509\,
            I => \N__12498\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__12506\,
            I => \N__12498\
        );

    \I__1444\ : LocalMux
    port map (
            O => \N__12503\,
            I => \uu0.l_precountZ0Z_0\
        );

    \I__1443\ : Odrv4
    port map (
            O => \N__12498\,
            I => \uu0.l_precountZ0Z_0\
        );

    \I__1442\ : InMux
    port map (
            O => \N__12493\,
            I => \N__12490\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__12490\,
            I => \N__12487\
        );

    \I__1440\ : Span4Mux_s1_v
    port map (
            O => \N__12487\,
            I => \N__12484\
        );

    \I__1439\ : Odrv4
    port map (
            O => \N__12484\,
            I => \uu0.un99_ci_0\
        );

    \I__1438\ : InMux
    port map (
            O => \N__12481\,
            I => \N__12475\
        );

    \I__1437\ : InMux
    port map (
            O => \N__12480\,
            I => \N__12475\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__12475\,
            I => \N__12470\
        );

    \I__1435\ : InMux
    port map (
            O => \N__12474\,
            I => \N__12467\
        );

    \I__1434\ : InMux
    port map (
            O => \N__12473\,
            I => \N__12464\
        );

    \I__1433\ : Span4Mux_h
    port map (
            O => \N__12470\,
            I => \N__12461\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__12467\,
            I => \N__12458\
        );

    \I__1431\ : LocalMux
    port map (
            O => \N__12464\,
            I => \uu0.l_countZ0Z_4\
        );

    \I__1430\ : Odrv4
    port map (
            O => \N__12461\,
            I => \uu0.l_countZ0Z_4\
        );

    \I__1429\ : Odrv4
    port map (
            O => \N__12458\,
            I => \uu0.l_countZ0Z_4\
        );

    \I__1428\ : InMux
    port map (
            O => \N__12451\,
            I => \N__12446\
        );

    \I__1427\ : InMux
    port map (
            O => \N__12450\,
            I => \N__12441\
        );

    \I__1426\ : InMux
    port map (
            O => \N__12449\,
            I => \N__12441\
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__12446\,
            I => \N__12438\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__12441\,
            I => \uu0.l_countZ0Z_5\
        );

    \I__1423\ : Odrv4
    port map (
            O => \N__12438\,
            I => \uu0.l_countZ0Z_5\
        );

    \I__1422\ : CascadeMux
    port map (
            O => \N__12433\,
            I => \N__12430\
        );

    \I__1421\ : InMux
    port map (
            O => \N__12430\,
            I => \N__12427\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__12427\,
            I => \N__12423\
        );

    \I__1419\ : InMux
    port map (
            O => \N__12426\,
            I => \N__12420\
        );

    \I__1418\ : Span4Mux_h
    port map (
            O => \N__12423\,
            I => \N__12417\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__12420\,
            I => \uu0.un88_ci_3\
        );

    \I__1416\ : Odrv4
    port map (
            O => \N__12417\,
            I => \uu0.un88_ci_3\
        );

    \I__1415\ : InMux
    port map (
            O => \N__12412\,
            I => \N__12406\
        );

    \I__1414\ : InMux
    port map (
            O => \N__12411\,
            I => \N__12406\
        );

    \I__1413\ : LocalMux
    port map (
            O => \N__12406\,
            I => \N__12403\
        );

    \I__1412\ : Span4Mux_v
    port map (
            O => \N__12403\,
            I => \N__12397\
        );

    \I__1411\ : InMux
    port map (
            O => \N__12402\,
            I => \N__12394\
        );

    \I__1410\ : InMux
    port map (
            O => \N__12401\,
            I => \N__12389\
        );

    \I__1409\ : InMux
    port map (
            O => \N__12400\,
            I => \N__12389\
        );

    \I__1408\ : Odrv4
    port map (
            O => \N__12397\,
            I => \uu0.un66_ci\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__12394\,
            I => \uu0.un66_ci\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__12389\,
            I => \uu0.un66_ci\
        );

    \I__1405\ : CascadeMux
    port map (
            O => \N__12382\,
            I => \uu0.un88_ci_3_cascade_\
        );

    \I__1404\ : InMux
    port map (
            O => \N__12379\,
            I => \N__12376\
        );

    \I__1403\ : LocalMux
    port map (
            O => \N__12376\,
            I => \N__12370\
        );

    \I__1402\ : InMux
    port map (
            O => \N__12375\,
            I => \N__12367\
        );

    \I__1401\ : InMux
    port map (
            O => \N__12374\,
            I => \N__12364\
        );

    \I__1400\ : InMux
    port map (
            O => \N__12373\,
            I => \N__12361\
        );

    \I__1399\ : Span4Mux_s3_h
    port map (
            O => \N__12370\,
            I => \N__12358\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__12367\,
            I => \N__12355\
        );

    \I__1397\ : LocalMux
    port map (
            O => \N__12364\,
            I => \uu0.l_countZ0Z_6\
        );

    \I__1396\ : LocalMux
    port map (
            O => \N__12361\,
            I => \uu0.l_countZ0Z_6\
        );

    \I__1395\ : Odrv4
    port map (
            O => \N__12358\,
            I => \uu0.l_countZ0Z_6\
        );

    \I__1394\ : Odrv4
    port map (
            O => \N__12355\,
            I => \uu0.l_countZ0Z_6\
        );

    \I__1393\ : CEMux
    port map (
            O => \N__12346\,
            I => \N__12331\
        );

    \I__1392\ : CEMux
    port map (
            O => \N__12345\,
            I => \N__12331\
        );

    \I__1391\ : CEMux
    port map (
            O => \N__12344\,
            I => \N__12331\
        );

    \I__1390\ : CEMux
    port map (
            O => \N__12343\,
            I => \N__12331\
        );

    \I__1389\ : CEMux
    port map (
            O => \N__12342\,
            I => \N__12331\
        );

    \I__1388\ : GlobalMux
    port map (
            O => \N__12331\,
            I => \N__12328\
        );

    \I__1387\ : gio2CtrlBuf
    port map (
            O => \N__12328\,
            I => \uu0.un11_l_count_i_g\
        );

    \I__1386\ : InMux
    port map (
            O => \N__12325\,
            I => \N__12322\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__12322\,
            I => \Lab_UT.dictrl.N_5_0_0\
        );

    \I__1384\ : CascadeMux
    port map (
            O => \N__12319\,
            I => \Lab_UT.dictrl.g0_4_0_cascade_\
        );

    \I__1383\ : CascadeMux
    port map (
            O => \N__12316\,
            I => \Lab_UT.dictrl.N_8_0_0_cascade_\
        );

    \I__1382\ : InMux
    port map (
            O => \N__12313\,
            I => \N__12310\
        );

    \I__1381\ : LocalMux
    port map (
            O => \N__12310\,
            I => \Lab_UT.dictrl.N_4\
        );

    \I__1380\ : InMux
    port map (
            O => \N__12307\,
            I => \N__12304\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__12304\,
            I => \Lab_UT.dictrl.currState_i_5_2\
        );

    \I__1378\ : CascadeMux
    port map (
            O => \N__12301\,
            I => \Lab_UT.dictrl.G_19_0_a7_4_10_cascade_\
        );

    \I__1377\ : CascadeMux
    port map (
            O => \N__12298\,
            I => \Lab_UT.dictrl.N_21_cascade_\
        );

    \I__1376\ : InMux
    port map (
            O => \N__12295\,
            I => \N__12292\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__12292\,
            I => \N__12289\
        );

    \I__1374\ : Odrv12
    port map (
            O => \N__12289\,
            I => \Lab_UT.dictrl.G_19_0_a7_2_0\
        );

    \I__1373\ : InMux
    port map (
            O => \N__12286\,
            I => \N__12283\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__12283\,
            I => \Lab_UT.dictrl.G_19_0_0\
        );

    \I__1371\ : CascadeMux
    port map (
            O => \N__12280\,
            I => \Lab_UT.dictrl.i8_mux_0_0_cascade_\
        );

    \I__1370\ : InMux
    port map (
            O => \N__12277\,
            I => \N__12274\
        );

    \I__1369\ : LocalMux
    port map (
            O => \N__12274\,
            I => \Lab_UT.dictrl.i7_mux_0\
        );

    \I__1368\ : InMux
    port map (
            O => \N__12271\,
            I => \N__12268\
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__12268\,
            I => \Lab_UT.dictrl.N_12\
        );

    \I__1366\ : InMux
    port map (
            O => \N__12265\,
            I => \N__12262\
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__12262\,
            I => \N__12259\
        );

    \I__1364\ : Odrv4
    port map (
            O => \N__12259\,
            I => \Lab_UT.dictrl.G_30_0_a7_2\
        );

    \I__1363\ : CascadeMux
    port map (
            O => \N__12256\,
            I => \Lab_UT.dictrl.N_11_0_cascade_\
        );

    \I__1362\ : CascadeMux
    port map (
            O => \N__12253\,
            I => \N__12250\
        );

    \I__1361\ : InMux
    port map (
            O => \N__12250\,
            I => \N__12247\
        );

    \I__1360\ : LocalMux
    port map (
            O => \N__12247\,
            I => \Lab_UT.dictrl.G_30_0_a7_4_1\
        );

    \I__1359\ : InMux
    port map (
            O => \N__12244\,
            I => \N__12241\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__12241\,
            I => \Lab_UT.dictrl.G_30_0_a7_1_2\
        );

    \I__1357\ : CascadeMux
    port map (
            O => \N__12238\,
            I => \Lab_UT.dictrl.N_31_0_cascade_\
        );

    \I__1356\ : InMux
    port map (
            O => \N__12235\,
            I => \N__12232\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__12232\,
            I => \Lab_UT.dictrl.N_23_1\
        );

    \I__1354\ : CascadeMux
    port map (
            O => \N__12229\,
            I => \Lab_UT.dictrl.G_30_0_2_cascade_\
        );

    \I__1353\ : CascadeMux
    port map (
            O => \N__12226\,
            I => \Lab_UT.dictrl.nextStateZ0Z_1_cascade_\
        );

    \I__1352\ : CascadeMux
    port map (
            O => \N__12223\,
            I => \Lab_UT.dictrl.G_30_0_a7_2_0_cascade_\
        );

    \I__1351\ : InMux
    port map (
            O => \N__12220\,
            I => \N__12217\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__12217\,
            I => \Lab_UT.dictrl.G_30_0_0\
        );

    \I__1349\ : InMux
    port map (
            O => \N__12214\,
            I => \N__12211\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__12211\,
            I => \Lab_UT.dictrl.G_30_0_a7_0_0\
        );

    \I__1347\ : InMux
    port map (
            O => \N__12208\,
            I => \N__12205\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__12205\,
            I => \Lab_UT.dictrl.N_30_0\
        );

    \I__1345\ : InMux
    port map (
            O => \N__12202\,
            I => \N__12187\
        );

    \I__1344\ : InMux
    port map (
            O => \N__12201\,
            I => \N__12187\
        );

    \I__1343\ : InMux
    port map (
            O => \N__12200\,
            I => \N__12187\
        );

    \I__1342\ : InMux
    port map (
            O => \N__12199\,
            I => \N__12187\
        );

    \I__1341\ : InMux
    port map (
            O => \N__12198\,
            I => \N__12187\
        );

    \I__1340\ : LocalMux
    port map (
            O => \N__12187\,
            I => \uu2.l_countZ0Z_6\
        );

    \I__1339\ : CascadeMux
    port map (
            O => \N__12184\,
            I => \N__12178\
        );

    \I__1338\ : InMux
    port map (
            O => \N__12183\,
            I => \N__12172\
        );

    \I__1337\ : InMux
    port map (
            O => \N__12182\,
            I => \N__12172\
        );

    \I__1336\ : InMux
    port map (
            O => \N__12181\,
            I => \N__12165\
        );

    \I__1335\ : InMux
    port map (
            O => \N__12178\,
            I => \N__12165\
        );

    \I__1334\ : InMux
    port map (
            O => \N__12177\,
            I => \N__12165\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__12172\,
            I => \uu2.l_countZ0Z_4\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__12165\,
            I => \uu2.l_countZ0Z_4\
        );

    \I__1331\ : CascadeMux
    port map (
            O => \N__12160\,
            I => \N__12155\
        );

    \I__1330\ : InMux
    port map (
            O => \N__12159\,
            I => \N__12148\
        );

    \I__1329\ : InMux
    port map (
            O => \N__12158\,
            I => \N__12148\
        );

    \I__1328\ : InMux
    port map (
            O => \N__12155\,
            I => \N__12148\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__12148\,
            I => \uu2.l_countZ0Z_9\
        );

    \I__1326\ : InMux
    port map (
            O => \N__12145\,
            I => \N__12142\
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__12142\,
            I => \uu2.un1_l_count_2_2\
        );

    \I__1324\ : CascadeMux
    port map (
            O => \N__12139\,
            I => \Lab_UT.dictrl.N_8_1_cascade_\
        );

    \I__1323\ : CascadeMux
    port map (
            O => \N__12136\,
            I => \Lab_UT.dictrl.N_20_0_cascade_\
        );

    \I__1322\ : InMux
    port map (
            O => \N__12133\,
            I => \N__12130\
        );

    \I__1321\ : LocalMux
    port map (
            O => \N__12130\,
            I => \Lab_UT.dictrl.N_9_1\
        );

    \I__1320\ : InMux
    port map (
            O => \N__12127\,
            I => \N__12112\
        );

    \I__1319\ : InMux
    port map (
            O => \N__12126\,
            I => \N__12112\
        );

    \I__1318\ : InMux
    port map (
            O => \N__12125\,
            I => \N__12112\
        );

    \I__1317\ : InMux
    port map (
            O => \N__12124\,
            I => \N__12112\
        );

    \I__1316\ : InMux
    port map (
            O => \N__12123\,
            I => \N__12112\
        );

    \I__1315\ : LocalMux
    port map (
            O => \N__12112\,
            I => \uu2.l_countZ0Z_2\
        );

    \I__1314\ : InMux
    port map (
            O => \N__12109\,
            I => \N__12100\
        );

    \I__1313\ : InMux
    port map (
            O => \N__12108\,
            I => \N__12100\
        );

    \I__1312\ : InMux
    port map (
            O => \N__12107\,
            I => \N__12100\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__12100\,
            I => \uu2.l_countZ0Z_3\
        );

    \I__1310\ : CascadeMux
    port map (
            O => \N__12097\,
            I => \uu2.un306_ci_cascade_\
        );

    \I__1309\ : CascadeMux
    port map (
            O => \N__12094\,
            I => \uu2.un350_ci_cascade_\
        );

    \I__1308\ : InMux
    port map (
            O => \N__12091\,
            I => \N__12088\
        );

    \I__1307\ : LocalMux
    port map (
            O => \N__12088\,
            I => \uu2.un1_l_count_1_2_0\
        );

    \I__1306\ : InMux
    port map (
            O => \N__12085\,
            I => \N__12082\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__12082\,
            I => \uu2.un350_ci\
        );

    \I__1304\ : CascadeMux
    port map (
            O => \N__12079\,
            I => \N__12074\
        );

    \I__1303\ : InMux
    port map (
            O => \N__12078\,
            I => \N__12071\
        );

    \I__1302\ : InMux
    port map (
            O => \N__12077\,
            I => \N__12068\
        );

    \I__1301\ : InMux
    port map (
            O => \N__12074\,
            I => \N__12065\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__12071\,
            I => \uu2.l_countZ0Z_8\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__12068\,
            I => \uu2.l_countZ0Z_8\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__12065\,
            I => \uu2.l_countZ0Z_8\
        );

    \I__1297\ : InMux
    port map (
            O => \N__12058\,
            I => \N__12053\
        );

    \I__1296\ : InMux
    port map (
            O => \N__12057\,
            I => \N__12048\
        );

    \I__1295\ : InMux
    port map (
            O => \N__12056\,
            I => \N__12048\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__12053\,
            I => \uu2.l_countZ0Z_5\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__12048\,
            I => \uu2.l_countZ0Z_5\
        );

    \I__1292\ : CascadeMux
    port map (
            O => \N__12043\,
            I => \N__12039\
        );

    \I__1291\ : CascadeMux
    port map (
            O => \N__12042\,
            I => \N__12036\
        );

    \I__1290\ : InMux
    port map (
            O => \N__12039\,
            I => \N__12031\
        );

    \I__1289\ : InMux
    port map (
            O => \N__12036\,
            I => \N__12031\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__12031\,
            I => \uu2.vbuf_count.un328_ci_3\
        );

    \I__1287\ : CascadeMux
    port map (
            O => \N__12028\,
            I => \uu2.vbuf_count.un328_ci_3_cascade_\
        );

    \I__1286\ : InMux
    port map (
            O => \N__12025\,
            I => \N__12019\
        );

    \I__1285\ : InMux
    port map (
            O => \N__12024\,
            I => \N__12012\
        );

    \I__1284\ : InMux
    port map (
            O => \N__12023\,
            I => \N__12012\
        );

    \I__1283\ : InMux
    port map (
            O => \N__12022\,
            I => \N__12012\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__12019\,
            I => \uu2.un306_ci\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__12012\,
            I => \uu2.un306_ci\
        );

    \I__1280\ : InMux
    port map (
            O => \N__12007\,
            I => \N__12000\
        );

    \I__1279\ : InMux
    port map (
            O => \N__12006\,
            I => \N__12000\
        );

    \I__1278\ : InMux
    port map (
            O => \N__12005\,
            I => \N__11997\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__12000\,
            I => \uu2.l_countZ0Z_7\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__11997\,
            I => \uu2.l_countZ0Z_7\
        );

    \I__1275\ : InMux
    port map (
            O => \N__11992\,
            I => \N__11989\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__11989\,
            I => vbuf_tx_data_4
        );

    \I__1273\ : InMux
    port map (
            O => \N__11986\,
            I => \N__11983\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__11983\,
            I => \buart.Z_tx.shifterZ0Z_5\
        );

    \I__1271\ : InMux
    port map (
            O => \N__11980\,
            I => \N__11977\
        );

    \I__1270\ : LocalMux
    port map (
            O => \N__11977\,
            I => vbuf_tx_data_5
        );

    \I__1269\ : InMux
    port map (
            O => \N__11974\,
            I => \N__11971\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__11971\,
            I => \buart.Z_tx.shifterZ0Z_6\
        );

    \I__1267\ : CascadeMux
    port map (
            O => \N__11968\,
            I => \uu2.un1_l_count_1_3_cascade_\
        );

    \I__1266\ : CascadeMux
    port map (
            O => \N__11965\,
            I => \N__11962\
        );

    \I__1265\ : InMux
    port map (
            O => \N__11962\,
            I => \N__11959\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__11959\,
            I => \uu2.un1_l_count_1_3\
        );

    \I__1263\ : CascadeMux
    port map (
            O => \N__11956\,
            I => \uu2.un1_l_count_2_0_cascade_\
        );

    \I__1262\ : InMux
    port map (
            O => \N__11953\,
            I => \N__11950\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__11950\,
            I => \uu2.r_data_wire_6\
        );

    \I__1260\ : InMux
    port map (
            O => \N__11947\,
            I => \N__11944\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__11944\,
            I => \uu2.r_data_wire_7\
        );

    \I__1258\ : InMux
    port map (
            O => \N__11941\,
            I => \N__11938\
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__11938\,
            I => vbuf_tx_data_0
        );

    \I__1256\ : InMux
    port map (
            O => \N__11935\,
            I => \N__11932\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__11932\,
            I => \buart.Z_tx.shifterZ0Z_1\
        );

    \I__1254\ : InMux
    port map (
            O => \N__11929\,
            I => \N__11926\
        );

    \I__1253\ : LocalMux
    port map (
            O => \N__11926\,
            I => \buart.Z_tx.shifterZ0Z_0\
        );

    \I__1252\ : IoInMux
    port map (
            O => \N__11923\,
            I => \N__11920\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__11920\,
            I => \N__11917\
        );

    \I__1250\ : Span4Mux_s1_h
    port map (
            O => \N__11917\,
            I => \N__11914\
        );

    \I__1249\ : Span4Mux_v
    port map (
            O => \N__11914\,
            I => \N__11911\
        );

    \I__1248\ : Odrv4
    port map (
            O => \N__11911\,
            I => o_serial_data_c
        );

    \I__1247\ : InMux
    port map (
            O => \N__11908\,
            I => \N__11905\
        );

    \I__1246\ : LocalMux
    port map (
            O => \N__11905\,
            I => vbuf_tx_data_1
        );

    \I__1245\ : InMux
    port map (
            O => \N__11902\,
            I => \N__11899\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__11899\,
            I => \buart.Z_tx.shifterZ0Z_2\
        );

    \I__1243\ : InMux
    port map (
            O => \N__11896\,
            I => \N__11893\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__11893\,
            I => vbuf_tx_data_2
        );

    \I__1241\ : InMux
    port map (
            O => \N__11890\,
            I => \N__11887\
        );

    \I__1240\ : LocalMux
    port map (
            O => \N__11887\,
            I => \buart.Z_tx.shifterZ0Z_3\
        );

    \I__1239\ : InMux
    port map (
            O => \N__11884\,
            I => \N__11881\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__11881\,
            I => vbuf_tx_data_3
        );

    \I__1237\ : InMux
    port map (
            O => \N__11878\,
            I => \N__11875\
        );

    \I__1236\ : LocalMux
    port map (
            O => \N__11875\,
            I => \buart.Z_tx.shifterZ0Z_4\
        );

    \I__1235\ : InMux
    port map (
            O => \N__11872\,
            I => \N__11857\
        );

    \I__1234\ : InMux
    port map (
            O => \N__11871\,
            I => \N__11857\
        );

    \I__1233\ : InMux
    port map (
            O => \N__11870\,
            I => \N__11857\
        );

    \I__1232\ : InMux
    port map (
            O => \N__11869\,
            I => \N__11857\
        );

    \I__1231\ : InMux
    port map (
            O => \N__11868\,
            I => \N__11857\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__11857\,
            I => \uu0.l_precountZ0Z_1\
        );

    \I__1229\ : CascadeMux
    port map (
            O => \N__11854\,
            I => \N__11849\
        );

    \I__1228\ : CascadeMux
    port map (
            O => \N__11853\,
            I => \N__11846\
        );

    \I__1227\ : InMux
    port map (
            O => \N__11852\,
            I => \N__11839\
        );

    \I__1226\ : InMux
    port map (
            O => \N__11849\,
            I => \N__11839\
        );

    \I__1225\ : InMux
    port map (
            O => \N__11846\,
            I => \N__11839\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__11839\,
            I => \uu0.l_precountZ0Z_3\
        );

    \I__1223\ : CascadeMux
    port map (
            O => \N__11836\,
            I => \N__11831\
        );

    \I__1222\ : InMux
    port map (
            O => \N__11835\,
            I => \N__11823\
        );

    \I__1221\ : InMux
    port map (
            O => \N__11834\,
            I => \N__11823\
        );

    \I__1220\ : InMux
    port map (
            O => \N__11831\,
            I => \N__11823\
        );

    \I__1219\ : InMux
    port map (
            O => \N__11830\,
            I => \N__11820\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__11823\,
            I => \uu0.l_countZ0Z_1\
        );

    \I__1217\ : LocalMux
    port map (
            O => \N__11820\,
            I => \uu0.l_countZ0Z_1\
        );

    \I__1216\ : InMux
    port map (
            O => \N__11815\,
            I => \N__11811\
        );

    \I__1215\ : InMux
    port map (
            O => \N__11814\,
            I => \N__11808\
        );

    \I__1214\ : LocalMux
    port map (
            O => \N__11811\,
            I => \uu0.l_countZ0Z_18\
        );

    \I__1213\ : LocalMux
    port map (
            O => \N__11808\,
            I => \uu0.l_countZ0Z_18\
        );

    \I__1212\ : InMux
    port map (
            O => \N__11803\,
            I => \N__11798\
        );

    \I__1211\ : InMux
    port map (
            O => \N__11802\,
            I => \N__11793\
        );

    \I__1210\ : InMux
    port map (
            O => \N__11801\,
            I => \N__11793\
        );

    \I__1209\ : LocalMux
    port map (
            O => \N__11798\,
            I => \N__11790\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__11793\,
            I => \uu0.l_countZ0Z_15\
        );

    \I__1207\ : Odrv4
    port map (
            O => \N__11790\,
            I => \uu0.l_countZ0Z_15\
        );

    \I__1206\ : CascadeMux
    port map (
            O => \N__11785\,
            I => \uu0.un4_l_count_11_cascade_\
        );

    \I__1205\ : InMux
    port map (
            O => \N__11782\,
            I => \N__11779\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__11779\,
            I => \N__11776\
        );

    \I__1203\ : Odrv4
    port map (
            O => \N__11776\,
            I => \uu0.un4_l_count_16\
        );

    \I__1202\ : InMux
    port map (
            O => \N__11773\,
            I => \N__11770\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__11770\,
            I => \uu2.r_data_wire_0\
        );

    \I__1200\ : InMux
    port map (
            O => \N__11767\,
            I => \N__11764\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__11764\,
            I => \uu2.r_data_wire_1\
        );

    \I__1198\ : InMux
    port map (
            O => \N__11761\,
            I => \N__11758\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__11758\,
            I => \uu2.r_data_wire_2\
        );

    \I__1196\ : InMux
    port map (
            O => \N__11755\,
            I => \N__11752\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__11752\,
            I => \uu2.r_data_wire_3\
        );

    \I__1194\ : InMux
    port map (
            O => \N__11749\,
            I => \N__11746\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__11746\,
            I => \uu2.r_data_wire_4\
        );

    \I__1192\ : InMux
    port map (
            O => \N__11743\,
            I => \N__11740\
        );

    \I__1191\ : LocalMux
    port map (
            O => \N__11740\,
            I => \uu2.r_data_wire_5\
        );

    \I__1190\ : CascadeMux
    port map (
            O => \N__11737\,
            I => \N__11729\
        );

    \I__1189\ : CascadeMux
    port map (
            O => \N__11736\,
            I => \N__11726\
        );

    \I__1188\ : CascadeMux
    port map (
            O => \N__11735\,
            I => \N__11720\
        );

    \I__1187\ : CascadeMux
    port map (
            O => \N__11734\,
            I => \N__11717\
        );

    \I__1186\ : InMux
    port map (
            O => \N__11733\,
            I => \N__11709\
        );

    \I__1185\ : InMux
    port map (
            O => \N__11732\,
            I => \N__11709\
        );

    \I__1184\ : InMux
    port map (
            O => \N__11729\,
            I => \N__11709\
        );

    \I__1183\ : InMux
    port map (
            O => \N__11726\,
            I => \N__11706\
        );

    \I__1182\ : InMux
    port map (
            O => \N__11725\,
            I => \N__11699\
        );

    \I__1181\ : InMux
    port map (
            O => \N__11724\,
            I => \N__11699\
        );

    \I__1180\ : InMux
    port map (
            O => \N__11723\,
            I => \N__11699\
        );

    \I__1179\ : InMux
    port map (
            O => \N__11720\,
            I => \N__11692\
        );

    \I__1178\ : InMux
    port map (
            O => \N__11717\,
            I => \N__11692\
        );

    \I__1177\ : InMux
    port map (
            O => \N__11716\,
            I => \N__11692\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__11709\,
            I => \uu0.un110_ci\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__11706\,
            I => \uu0.un110_ci\
        );

    \I__1174\ : LocalMux
    port map (
            O => \N__11699\,
            I => \uu0.un110_ci\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__11692\,
            I => \uu0.un110_ci\
        );

    \I__1172\ : InMux
    port map (
            O => \N__11683\,
            I => \N__11676\
        );

    \I__1171\ : InMux
    port map (
            O => \N__11682\,
            I => \N__11676\
        );

    \I__1170\ : InMux
    port map (
            O => \N__11681\,
            I => \N__11673\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__11676\,
            I => \N__11670\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__11673\,
            I => \uu0.un198_ci_2\
        );

    \I__1167\ : Odrv4
    port map (
            O => \N__11670\,
            I => \uu0.un198_ci_2\
        );

    \I__1166\ : CascadeMux
    port map (
            O => \N__11665\,
            I => \uu0.un110_ci_cascade_\
        );

    \I__1165\ : InMux
    port map (
            O => \N__11662\,
            I => \N__11654\
        );

    \I__1164\ : InMux
    port map (
            O => \N__11661\,
            I => \N__11654\
        );

    \I__1163\ : InMux
    port map (
            O => \N__11660\,
            I => \N__11649\
        );

    \I__1162\ : InMux
    port map (
            O => \N__11659\,
            I => \N__11649\
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__11654\,
            I => \uu0.l_countZ0Z_16\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__11649\,
            I => \uu0.l_countZ0Z_16\
        );

    \I__1159\ : CascadeMux
    port map (
            O => \N__11644\,
            I => \uu0.un220_ci_cascade_\
        );

    \I__1158\ : InMux
    port map (
            O => \N__11641\,
            I => \N__11630\
        );

    \I__1157\ : InMux
    port map (
            O => \N__11640\,
            I => \N__11630\
        );

    \I__1156\ : InMux
    port map (
            O => \N__11639\,
            I => \N__11630\
        );

    \I__1155\ : InMux
    port map (
            O => \N__11638\,
            I => \N__11625\
        );

    \I__1154\ : InMux
    port map (
            O => \N__11637\,
            I => \N__11625\
        );

    \I__1153\ : LocalMux
    port map (
            O => \N__11630\,
            I => \uu0.l_countZ0Z_9\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__11625\,
            I => \uu0.l_countZ0Z_9\
        );

    \I__1151\ : CascadeMux
    port map (
            O => \N__11620\,
            I => \N__11617\
        );

    \I__1150\ : InMux
    port map (
            O => \N__11617\,
            I => \N__11608\
        );

    \I__1149\ : InMux
    port map (
            O => \N__11616\,
            I => \N__11608\
        );

    \I__1148\ : InMux
    port map (
            O => \N__11615\,
            I => \N__11608\
        );

    \I__1147\ : LocalMux
    port map (
            O => \N__11608\,
            I => \uu0.l_countZ0Z_7\
        );

    \I__1146\ : CascadeMux
    port map (
            O => \N__11605\,
            I => \N__11600\
        );

    \I__1145\ : InMux
    port map (
            O => \N__11604\,
            I => \N__11593\
        );

    \I__1144\ : InMux
    port map (
            O => \N__11603\,
            I => \N__11593\
        );

    \I__1143\ : InMux
    port map (
            O => \N__11600\,
            I => \N__11593\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__11593\,
            I => \uu0.l_countZ0Z_17\
        );

    \I__1141\ : InMux
    port map (
            O => \N__11590\,
            I => \N__11583\
        );

    \I__1140\ : InMux
    port map (
            O => \N__11589\,
            I => \N__11583\
        );

    \I__1139\ : InMux
    port map (
            O => \N__11588\,
            I => \N__11580\
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__11583\,
            I => \uu0.l_countZ0Z_3\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__11580\,
            I => \uu0.l_countZ0Z_3\
        );

    \I__1136\ : InMux
    port map (
            O => \N__11575\,
            I => \N__11572\
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__11572\,
            I => \uu0.un4_l_count_12\
        );

    \I__1134\ : InMux
    port map (
            O => \N__11569\,
            I => \N__11566\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__11566\,
            I => \N__11560\
        );

    \I__1132\ : InMux
    port map (
            O => \N__11565\,
            I => \N__11557\
        );

    \I__1131\ : CascadeMux
    port map (
            O => \N__11564\,
            I => \N__11554\
        );

    \I__1130\ : CascadeMux
    port map (
            O => \N__11563\,
            I => \N__11551\
        );

    \I__1129\ : Span4Mux_s2_v
    port map (
            O => \N__11560\,
            I => \N__11547\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__11557\,
            I => \N__11544\
        );

    \I__1127\ : InMux
    port map (
            O => \N__11554\,
            I => \N__11537\
        );

    \I__1126\ : InMux
    port map (
            O => \N__11551\,
            I => \N__11537\
        );

    \I__1125\ : InMux
    port map (
            O => \N__11550\,
            I => \N__11537\
        );

    \I__1124\ : Odrv4
    port map (
            O => \N__11547\,
            I => \buart.Z_tx.uart_busy_0_i\
        );

    \I__1123\ : Odrv4
    port map (
            O => \N__11544\,
            I => \buart.Z_tx.uart_busy_0_i\
        );

    \I__1122\ : LocalMux
    port map (
            O => \N__11537\,
            I => \buart.Z_tx.uart_busy_0_i\
        );

    \I__1121\ : InMux
    port map (
            O => \N__11530\,
            I => \N__11527\
        );

    \I__1120\ : LocalMux
    port map (
            O => \N__11527\,
            I => \N__11520\
        );

    \I__1119\ : InMux
    port map (
            O => \N__11526\,
            I => \N__11513\
        );

    \I__1118\ : InMux
    port map (
            O => \N__11525\,
            I => \N__11506\
        );

    \I__1117\ : InMux
    port map (
            O => \N__11524\,
            I => \N__11506\
        );

    \I__1116\ : InMux
    port map (
            O => \N__11523\,
            I => \N__11506\
        );

    \I__1115\ : Span4Mux_s2_v
    port map (
            O => \N__11520\,
            I => \N__11503\
        );

    \I__1114\ : InMux
    port map (
            O => \N__11519\,
            I => \N__11494\
        );

    \I__1113\ : InMux
    port map (
            O => \N__11518\,
            I => \N__11494\
        );

    \I__1112\ : InMux
    port map (
            O => \N__11517\,
            I => \N__11494\
        );

    \I__1111\ : InMux
    port map (
            O => \N__11516\,
            I => \N__11494\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__11513\,
            I => \N__11491\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__11506\,
            I => \buart.Z_tx.ser_clk\
        );

    \I__1108\ : Odrv4
    port map (
            O => \N__11503\,
            I => \buart.Z_tx.ser_clk\
        );

    \I__1107\ : LocalMux
    port map (
            O => \N__11494\,
            I => \buart.Z_tx.ser_clk\
        );

    \I__1106\ : Odrv12
    port map (
            O => \N__11491\,
            I => \buart.Z_tx.ser_clk\
        );

    \I__1105\ : CascadeMux
    port map (
            O => \N__11482\,
            I => \N__11477\
        );

    \I__1104\ : InMux
    port map (
            O => \N__11481\,
            I => \N__11474\
        );

    \I__1103\ : InMux
    port map (
            O => \N__11480\,
            I => \N__11471\
        );

    \I__1102\ : InMux
    port map (
            O => \N__11477\,
            I => \N__11468\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__11474\,
            I => \N__11465\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__11471\,
            I => \buart.Z_tx.bitcountZ0Z_0\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__11468\,
            I => \buart.Z_tx.bitcountZ0Z_0\
        );

    \I__1098\ : Odrv4
    port map (
            O => \N__11465\,
            I => \buart.Z_tx.bitcountZ0Z_0\
        );

    \I__1097\ : CascadeMux
    port map (
            O => \N__11458\,
            I => \N__11452\
        );

    \I__1096\ : InMux
    port map (
            O => \N__11457\,
            I => \N__11445\
        );

    \I__1095\ : InMux
    port map (
            O => \N__11456\,
            I => \N__11445\
        );

    \I__1094\ : InMux
    port map (
            O => \N__11455\,
            I => \N__11445\
        );

    \I__1093\ : InMux
    port map (
            O => \N__11452\,
            I => \N__11442\
        );

    \I__1092\ : LocalMux
    port map (
            O => \N__11445\,
            I => \uu0.l_precountZ0Z_2\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__11442\,
            I => \uu0.l_precountZ0Z_2\
        );

    \I__1090\ : InMux
    port map (
            O => \N__11437\,
            I => \N__11434\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__11434\,
            I => \uu0.un4_l_count_13\
        );

    \I__1088\ : CascadeMux
    port map (
            O => \N__11431\,
            I => \uu0.un4_l_count_18_cascade_\
        );

    \I__1087\ : CascadeMux
    port map (
            O => \N__11428\,
            I => \uu0.un4_l_count_0_cascade_\
        );

    \I__1086\ : InMux
    port map (
            O => \N__11425\,
            I => \N__11422\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__11422\,
            I => \uu0.un143_ci_0\
        );

    \I__1084\ : CascadeMux
    port map (
            O => \N__11419\,
            I => \N__11415\
        );

    \I__1083\ : InMux
    port map (
            O => \N__11418\,
            I => \N__11409\
        );

    \I__1082\ : InMux
    port map (
            O => \N__11415\,
            I => \N__11409\
        );

    \I__1081\ : InMux
    port map (
            O => \N__11414\,
            I => \N__11406\
        );

    \I__1080\ : LocalMux
    port map (
            O => \N__11409\,
            I => \uu0.l_countZ0Z_11\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__11406\,
            I => \uu0.l_countZ0Z_11\
        );

    \I__1078\ : CascadeMux
    port map (
            O => \N__11401\,
            I => \N__11398\
        );

    \I__1077\ : InMux
    port map (
            O => \N__11398\,
            I => \N__11386\
        );

    \I__1076\ : InMux
    port map (
            O => \N__11397\,
            I => \N__11386\
        );

    \I__1075\ : InMux
    port map (
            O => \N__11396\,
            I => \N__11386\
        );

    \I__1074\ : InMux
    port map (
            O => \N__11395\,
            I => \N__11386\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__11386\,
            I => \uu0.l_countZ0Z_10\
        );

    \I__1072\ : InMux
    port map (
            O => \N__11383\,
            I => \N__11375\
        );

    \I__1071\ : InMux
    port map (
            O => \N__11382\,
            I => \N__11375\
        );

    \I__1070\ : InMux
    port map (
            O => \N__11381\,
            I => \N__11370\
        );

    \I__1069\ : InMux
    port map (
            O => \N__11380\,
            I => \N__11370\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__11375\,
            I => \uu0.un154_ci_9\
        );

    \I__1067\ : LocalMux
    port map (
            O => \N__11370\,
            I => \uu0.un154_ci_9\
        );

    \I__1066\ : CascadeMux
    port map (
            O => \N__11365\,
            I => \uu0.un154_ci_9_cascade_\
        );

    \I__1065\ : InMux
    port map (
            O => \N__11362\,
            I => \N__11357\
        );

    \I__1064\ : InMux
    port map (
            O => \N__11361\,
            I => \N__11352\
        );

    \I__1063\ : InMux
    port map (
            O => \N__11360\,
            I => \N__11352\
        );

    \I__1062\ : LocalMux
    port map (
            O => \N__11357\,
            I => \uu0.un4_l_count_0_8\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__11352\,
            I => \uu0.un4_l_count_0_8\
        );

    \I__1060\ : CascadeMux
    port map (
            O => \N__11347\,
            I => \N__11341\
        );

    \I__1059\ : InMux
    port map (
            O => \N__11346\,
            I => \N__11336\
        );

    \I__1058\ : InMux
    port map (
            O => \N__11345\,
            I => \N__11336\
        );

    \I__1057\ : InMux
    port map (
            O => \N__11344\,
            I => \N__11331\
        );

    \I__1056\ : InMux
    port map (
            O => \N__11341\,
            I => \N__11331\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__11336\,
            I => \uu0.l_countZ0Z_14\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__11331\,
            I => \uu0.l_countZ0Z_14\
        );

    \I__1053\ : InMux
    port map (
            O => \N__11326\,
            I => \N__11318\
        );

    \I__1052\ : InMux
    port map (
            O => \N__11325\,
            I => \N__11313\
        );

    \I__1051\ : InMux
    port map (
            O => \N__11324\,
            I => \N__11313\
        );

    \I__1050\ : InMux
    port map (
            O => \N__11323\,
            I => \N__11306\
        );

    \I__1049\ : InMux
    port map (
            O => \N__11322\,
            I => \N__11306\
        );

    \I__1048\ : InMux
    port map (
            O => \N__11321\,
            I => \N__11306\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__11318\,
            I => \uu0.l_countZ0Z_8\
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__11313\,
            I => \uu0.l_countZ0Z_8\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__11306\,
            I => \uu0.l_countZ0Z_8\
        );

    \I__1044\ : CascadeMux
    port map (
            O => \N__11299\,
            I => \Lab_UT.dictrl.currState_0_ret_28_RNOZ0Z_4_cascade_\
        );

    \I__1043\ : InMux
    port map (
            O => \N__11296\,
            I => \N__11293\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__11293\,
            I => \Lab_UT.dictrl.N_1605_0\
        );

    \I__1041\ : InMux
    port map (
            O => \N__11290\,
            I => \N__11287\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__11287\,
            I => \Lab_UT.dictrl.N_5_0\
        );

    \I__1039\ : CascadeMux
    port map (
            O => \N__11284\,
            I => \Lab_UT.dictrl.g1_0_cascade_\
        );

    \I__1038\ : CascadeMux
    port map (
            O => \N__11281\,
            I => \Lab_UT.dictrl.g0_i_o4_4_1_cascade_\
        );

    \I__1037\ : CascadeMux
    port map (
            O => \N__11278\,
            I => \Lab_UT.dictrl.g0_i_o4_4_cascade_\
        );

    \I__1036\ : InMux
    port map (
            O => \N__11275\,
            I => \N__11272\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__11272\,
            I => \uart_RXD\
        );

    \I__1034\ : InMux
    port map (
            O => \N__11269\,
            I => \N__11259\
        );

    \I__1033\ : InMux
    port map (
            O => \N__11268\,
            I => \N__11259\
        );

    \I__1032\ : InMux
    port map (
            O => \N__11267\,
            I => \N__11259\
        );

    \I__1031\ : InMux
    port map (
            O => \N__11266\,
            I => \N__11256\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__11259\,
            I => \uu0.l_countZ0Z_2\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__11256\,
            I => \uu0.l_countZ0Z_2\
        );

    \I__1028\ : CascadeMux
    port map (
            O => \N__11251\,
            I => \uu0.un4_l_count_14_cascade_\
        );

    \I__1027\ : CascadeMux
    port map (
            O => \N__11248\,
            I => \Lab_UT.dictrl.N_17_1_cascade_\
        );

    \I__1026\ : CascadeMux
    port map (
            O => \N__11245\,
            I => \Lab_UT.dictrl.g0_i_4_0_cascade_\
        );

    \I__1025\ : InMux
    port map (
            O => \N__11242\,
            I => \N__11239\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__11239\,
            I => \Lab_UT.dictrl.N_19\
        );

    \I__1023\ : CascadeMux
    port map (
            O => \N__11236\,
            I => \N__11233\
        );

    \I__1022\ : InMux
    port map (
            O => \N__11233\,
            I => \N__11230\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__11230\,
            I => \Lab_UT.dictrl.N_8_2\
        );

    \I__1020\ : CascadeMux
    port map (
            O => \N__11227\,
            I => \Lab_UT.dictrl.N_8_2_cascade_\
        );

    \I__1019\ : InMux
    port map (
            O => \N__11224\,
            I => \N__11221\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__11221\,
            I => \Lab_UT.dictrl.g0_i_a8_0_1\
        );

    \I__1017\ : InMux
    port map (
            O => \N__11218\,
            I => \N__11215\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__11215\,
            I => \Lab_UT.dictrl.N_1605_1\
        );

    \I__1015\ : InMux
    port map (
            O => \N__11212\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_2\
        );

    \I__1014\ : InMux
    port map (
            O => \N__11209\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_3\
        );

    \I__1013\ : InMux
    port map (
            O => \N__11206\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_4\
        );

    \I__1012\ : InMux
    port map (
            O => \N__11203\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_5\
        );

    \I__1011\ : CascadeMux
    port map (
            O => \N__11200\,
            I => \N__11197\
        );

    \I__1010\ : InMux
    port map (
            O => \N__11197\,
            I => \N__11191\
        );

    \I__1009\ : InMux
    port map (
            O => \N__11196\,
            I => \N__11191\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__11191\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_5\
        );

    \I__1007\ : CascadeMux
    port map (
            O => \N__11188\,
            I => \N__11185\
        );

    \I__1006\ : InMux
    port map (
            O => \N__11185\,
            I => \N__11179\
        );

    \I__1005\ : InMux
    port map (
            O => \N__11184\,
            I => \N__11179\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__11179\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_4\
        );

    \I__1003\ : CascadeMux
    port map (
            O => \N__11176\,
            I => \N__11172\
        );

    \I__1002\ : InMux
    port map (
            O => \N__11175\,
            I => \N__11169\
        );

    \I__1001\ : InMux
    port map (
            O => \N__11172\,
            I => \N__11166\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__11169\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_6\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__11166\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_6\
        );

    \I__998\ : InMux
    port map (
            O => \N__11161\,
            I => \N__11155\
        );

    \I__997\ : InMux
    port map (
            O => \N__11160\,
            I => \N__11155\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__11155\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_3\
        );

    \I__995\ : InMux
    port map (
            O => \N__11152\,
            I => \N__11146\
        );

    \I__994\ : InMux
    port map (
            O => \N__11151\,
            I => \N__11146\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__11146\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_2\
        );

    \I__992\ : CascadeMux
    port map (
            O => \N__11143\,
            I => \buart.Z_tx.Z_baudgen.ser_clk_4_cascade_\
        );

    \I__991\ : CascadeMux
    port map (
            O => \N__11140\,
            I => \N__11136\
        );

    \I__990\ : InMux
    port map (
            O => \N__11139\,
            I => \N__11132\
        );

    \I__989\ : InMux
    port map (
            O => \N__11136\,
            I => \N__11127\
        );

    \I__988\ : InMux
    port map (
            O => \N__11135\,
            I => \N__11127\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__11132\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_1\
        );

    \I__986\ : LocalMux
    port map (
            O => \N__11127\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_1\
        );

    \I__985\ : InMux
    port map (
            O => \N__11122\,
            I => \N__11114\
        );

    \I__984\ : InMux
    port map (
            O => \N__11121\,
            I => \N__11114\
        );

    \I__983\ : InMux
    port map (
            O => \N__11120\,
            I => \N__11109\
        );

    \I__982\ : InMux
    port map (
            O => \N__11119\,
            I => \N__11109\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__11114\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_0\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__11109\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_0\
        );

    \I__979\ : InMux
    port map (
            O => \N__11104\,
            I => \buart.Z_tx.un1_bitcount_cry_1\
        );

    \I__978\ : InMux
    port map (
            O => \N__11101\,
            I => \buart.Z_tx.un1_bitcount_cry_2\
        );

    \I__977\ : InMux
    port map (
            O => \N__11098\,
            I => \N__11095\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__11095\,
            I => \buart.Z_tx.bitcount_RNIVE1P1Z0Z_3\
        );

    \I__975\ : InMux
    port map (
            O => \N__11092\,
            I => \N__11089\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__11089\,
            I => \buart.Z_tx.un1_bitcount_axb_3\
        );

    \I__973\ : InMux
    port map (
            O => \N__11086\,
            I => \N__11083\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__11083\,
            I => \buart.Z_tx.un1_bitcount_cry_0_0_c_RNOZ0\
        );

    \I__971\ : CascadeMux
    port map (
            O => \N__11080\,
            I => \N__11077\
        );

    \I__970\ : InMux
    port map (
            O => \N__11077\,
            I => \N__11073\
        );

    \I__969\ : InMux
    port map (
            O => \N__11076\,
            I => \N__11070\
        );

    \I__968\ : LocalMux
    port map (
            O => \N__11073\,
            I => \buart.Z_tx.bitcountZ0Z_1\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__11070\,
            I => \buart.Z_tx.bitcountZ0Z_1\
        );

    \I__966\ : CascadeMux
    port map (
            O => \N__11065\,
            I => \N__11061\
        );

    \I__965\ : InMux
    port map (
            O => \N__11064\,
            I => \N__11058\
        );

    \I__964\ : InMux
    port map (
            O => \N__11061\,
            I => \N__11055\
        );

    \I__963\ : LocalMux
    port map (
            O => \N__11058\,
            I => \buart.Z_tx.bitcountZ0Z_3\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__11055\,
            I => \buart.Z_tx.bitcountZ0Z_3\
        );

    \I__961\ : CascadeMux
    port map (
            O => \N__11050\,
            I => \N__11047\
        );

    \I__960\ : InMux
    port map (
            O => \N__11047\,
            I => \N__11043\
        );

    \I__959\ : InMux
    port map (
            O => \N__11046\,
            I => \N__11040\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__11043\,
            I => \buart.Z_tx.bitcountZ0Z_2\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__11040\,
            I => \buart.Z_tx.bitcountZ0Z_2\
        );

    \I__956\ : CascadeMux
    port map (
            O => \N__11035\,
            I => \buart.Z_tx.uart_busy_0_i_cascade_\
        );

    \I__955\ : InMux
    port map (
            O => \N__11032\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_1\
        );

    \I__954\ : CascadeMux
    port map (
            O => \N__11029\,
            I => \N__11024\
        );

    \I__953\ : InMux
    port map (
            O => \N__11028\,
            I => \N__11011\
        );

    \I__952\ : InMux
    port map (
            O => \N__11027\,
            I => \N__11011\
        );

    \I__951\ : InMux
    port map (
            O => \N__11024\,
            I => \N__11011\
        );

    \I__950\ : InMux
    port map (
            O => \N__11023\,
            I => \N__11011\
        );

    \I__949\ : InMux
    port map (
            O => \N__11022\,
            I => \N__11011\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__11011\,
            I => \uu0.l_countZ0Z_0\
        );

    \I__947\ : CascadeMux
    port map (
            O => \N__11008\,
            I => \N__11005\
        );

    \I__946\ : InMux
    port map (
            O => \N__11005\,
            I => \N__11002\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__11002\,
            I => \uu0.un44_ci\
        );

    \I__944\ : CascadeMux
    port map (
            O => \N__10999\,
            I => \uu0.un44_ci_cascade_\
        );

    \I__943\ : InMux
    port map (
            O => \N__10996\,
            I => \buart.Z_tx.un1_bitcount_cry_0\
        );

    \I__942\ : InMux
    port map (
            O => \N__10993\,
            I => \N__10990\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__10990\,
            I => \buart.Z_tx.bitcount_RNIVE1P1_0Z0Z_3\
        );

    \I__940\ : CascadeMux
    port map (
            O => \N__10987\,
            I => \uu0.un187_ci_1_cascade_\
        );

    \I__939\ : InMux
    port map (
            O => \N__10984\,
            I => \N__10981\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__10981\,
            I => \uu0.un165_ci_0\
        );

    \I__937\ : CascadeMux
    port map (
            O => \N__10978\,
            I => \N__10975\
        );

    \I__936\ : InMux
    port map (
            O => \N__10975\,
            I => \N__10969\
        );

    \I__935\ : InMux
    port map (
            O => \N__10974\,
            I => \N__10969\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__10969\,
            I => \uu0.l_countZ0Z_13\
        );

    \I__933\ : InMux
    port map (
            O => \N__10966\,
            I => \N__10957\
        );

    \I__932\ : InMux
    port map (
            O => \N__10965\,
            I => \N__10957\
        );

    \I__931\ : InMux
    port map (
            O => \N__10964\,
            I => \N__10957\
        );

    \I__930\ : LocalMux
    port map (
            O => \N__10957\,
            I => \uu0.l_countZ0Z_12\
        );

    \I__929\ : CascadeMux
    port map (
            O => \N__10954\,
            I => \uu0.un4_l_count_0_8_cascade_\
        );

    \I__928\ : IoInMux
    port map (
            O => \N__10951\,
            I => \N__10948\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__10948\,
            I => \N__10945\
        );

    \I__926\ : Span12Mux_s9_v
    port map (
            O => \N__10945\,
            I => \N__10942\
        );

    \I__925\ : Odrv12
    port map (
            O => \N__10942\,
            I => \latticehx1k_pll_inst.clk\
        );

    \I__924\ : IoInMux
    port map (
            O => \N__10939\,
            I => \N__10936\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__10936\,
            I => \N__10933\
        );

    \I__922\ : IoSpan4Mux
    port map (
            O => \N__10933\,
            I => \N__10930\
        );

    \I__921\ : Odrv4
    port map (
            O => \N__10930\,
            I => clk_in_c
        );

    \INVuu2.w_addr_user_5C\ : INV
    port map (
            O => \INVuu2.w_addr_user_5C_net\,
            I => \N__29465\
        );

    \INVuu2.bitmap_93C\ : INV
    port map (
            O => \INVuu2.bitmap_93C_net\,
            I => \N__29435\
        );

    \INVuu2.w_addr_user_0C\ : INV
    port map (
            O => \INVuu2.w_addr_user_0C_net\,
            I => \N__29449\
        );

    \INVuu2.bitmap_212C\ : INV
    port map (
            O => \INVuu2.bitmap_212C_net\,
            I => \N__29416\
        );

    \INVuu2.bitmap_90C\ : INV
    port map (
            O => \INVuu2.bitmap_90C_net\,
            I => \N__29425\
        );

    \INVuu2.bitmap_308C\ : INV
    port map (
            O => \INVuu2.bitmap_308C_net\,
            I => \N__29434\
        );

    \INVuu2.w_addr_displaying_8C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_8C_net\,
            I => \N__29440\
        );

    \INVuu2.w_addr_user_nesr_3C\ : INV
    port map (
            O => \INVuu2.w_addr_user_nesr_3C_net\,
            I => \N__29448\
        );

    \INVuu2.bitmap_194C\ : INV
    port map (
            O => \INVuu2.bitmap_194C_net\,
            I => \N__29398\
        );

    \INVuu2.bitmap_203C\ : INV
    port map (
            O => \INVuu2.bitmap_203C_net\,
            I => \N__29404\
        );

    \INVuu2.bitmap_87C\ : INV
    port map (
            O => \INVuu2.bitmap_87C_net\,
            I => \N__29411\
        );

    \INVuu2.w_addr_displaying_nesr_3C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_nesr_3C_net\,
            I => \N__29418\
        );

    \INVuu2.bitmap_111C\ : INV
    port map (
            O => \INVuu2.bitmap_111C_net\,
            I => \N__29428\
        );

    \INVuu2.bitmap_72C\ : INV
    port map (
            O => \INVuu2.bitmap_72C_net\,
            I => \N__29415\
        );

    \INVuu2.bitmap_197C\ : INV
    port map (
            O => \INVuu2.bitmap_197C_net\,
            I => \N__29424\
        );

    \INVuu2.bitmap_290C\ : INV
    port map (
            O => \INVuu2.bitmap_290C_net\,
            I => \N__29433\
        );

    \INVuu2.vram_rd_clk_det_0C\ : INV
    port map (
            O => \INVuu2.vram_rd_clk_det_0C_net\,
            I => \N__29446\
        );

    \INVuu2.r_data_reg_0C\ : INV
    port map (
            O => \INVuu2.r_data_reg_0C_net\,
            I => \N__29460\
        );

    \IN_MUX_bfv_1_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_4_0_\
        );

    \IN_MUX_bfv_1_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_6_0_\
        );

    \IN_MUX_bfv_6_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_16_0_\
        );

    \IN_MUX_bfv_4_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_16_0_\
        );

    \IN_MUX_bfv_12_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_9_0_\
        );

    \latticehx1k_pll_inst.latticehx1k_pll_inst_RNIQV8B\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__10951\,
            GLOBALBUFFEROUTPUT => clk_g
        );

    \buart.Z_rx.bitcount_es_RNIV4M42_0_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__15649\,
            GLOBALBUFFEROUTPUT => \buart.Z_rx.sample_g\
        );

    \Lab_UT.uu0.delay_line_RNII8EF5_0_1\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__19111\,
            GLOBALBUFFEROUTPUT => \Lab_UT.uu0.un11_l_count_i_g\
        );

    \uu0.delay_line_RNILLLG7_0_1\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__12712\,
            GLOBALBUFFEROUTPUT => \uu0.un11_l_count_i_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \resetGen.rst_RNI4PQ1\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__24702\,
            GLOBALBUFFEROUTPUT => rst_g
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \uu0.l_count_13_LC_1_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001010001010000"
        )
    port map (
            in0 => \N__12982\,
            in1 => \N__10984\,
            in2 => \N__10978\,
            in3 => \N__11732\,
            lcout => \uu0.l_countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29480\,
            ce => \N__12343\,
            sr => \N__26085\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_1_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__11346\,
            in1 => \N__11381\,
            in2 => \_gnd_net_\,
            in3 => \N__11362\,
            lcout => OPEN,
            ltout => \uu0.un187_ci_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_15_LC_1_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001010101000000"
        )
    port map (
            in0 => \N__12983\,
            in1 => \N__11733\,
            in2 => \N__10987\,
            in3 => \N__11802\,
            lcout => \uu0.l_countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29480\,
            ce => \N__12343\,
            sr => \N__26085\
        );

    \uu0.l_count_12_LC_1_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__11383\,
            in1 => \N__10966\,
            in2 => \N__11737\,
            in3 => \N__12981\,
            lcout => \uu0.l_countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29480\,
            ce => \N__12343\,
            sr => \N__26085\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_1_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10965\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11382\,
            lcout => \uu0.un165_ci_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_RNIFAQ9_13_LC_1_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10974\,
            in2 => \_gnd_net_\,
            in3 => \N__10964\,
            lcout => \uu0.un4_l_count_0_8\,
            ltout => \uu0.un4_l_count_0_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_1_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__11380\,
            in1 => \N__11801\,
            in2 => \N__10954\,
            in3 => \N__11345\,
            lcout => \uu0.un198_ci_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_4_LC_1_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__12402\,
            in1 => \N__12473\,
            in2 => \_gnd_net_\,
            in3 => \N__12984\,
            lcout => \uu0.l_countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29480\,
            ce => \N__12343\,
            sr => \N__26085\
        );

    \uu0.l_count_RNI2CNU_11_LC_1_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__11414\,
            in1 => \N__11659\,
            in2 => \N__11458\,
            in3 => \N__11022\,
            lcout => \uu0.un4_l_count_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_3_LC_1_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__11269\,
            in1 => \N__11590\,
            in2 => \N__11008\,
            in3 => \N__12989\,
            lcout => \uu0.l_countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29478\,
            ce => \N__12342\,
            sr => \N__26083\
        );

    \uu0.l_count_1_LC_1_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__11835\,
            in1 => \N__11028\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uu0.l_countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29478\,
            ce => \N__12342\,
            sr => \N__26083\
        );

    \uu0.l_count_0_LC_1_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__11027\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12987\,
            lcout => \uu0.l_countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29478\,
            ce => \N__12342\,
            sr => \N__26083\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_1_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__11589\,
            in1 => \N__11267\,
            in2 => \N__11836\,
            in3 => \N__11023\,
            lcout => \uu0.un66_ci\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_1_LC_1_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11029\,
            in3 => \N__11834\,
            lcout => \uu0.un44_ci\,
            ltout => \uu0.un44_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_2_LC_1_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10999\,
            in3 => \N__11268\,
            lcout => \uu0.l_countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29478\,
            ce => \N__12342\,
            sr => \N__26083\
        );

    \uu0.l_count_16_LC_1_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__11660\,
            in1 => \N__11681\,
            in2 => \N__11736\,
            in3 => \N__12988\,
            lcout => \uu0.l_countZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29478\,
            ce => \N__12342\,
            sr => \N__26083\
        );

    \buart.Z_tx.bitcount_RNIVE1P1_0_3_LC_1_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11565\,
            in2 => \_gnd_net_\,
            in3 => \N__11526\,
            lcout => \buart.Z_tx.bitcount_RNIVE1P1_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.un1_bitcount_cry_0_0_c_LC_1_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11086\,
            in2 => \N__11482\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_4_0_\,
            carryout => \buart.Z_tx.un1_bitcount_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_1_LC_1_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__12825\,
            in1 => \N__11098\,
            in2 => \N__11080\,
            in3 => \N__10996\,
            lcout => \buart.Z_tx.bitcountZ0Z_1\,
            ltout => OPEN,
            carryin => \buart.Z_tx.un1_bitcount_cry_0\,
            carryout => \buart.Z_tx.un1_bitcount_cry_1\,
            clk => \N__29468\,
            ce => 'H',
            sr => \N__26079\
        );

    \buart.Z_tx.bitcount_2_LC_1_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__12811\,
            in1 => \N__10993\,
            in2 => \N__11050\,
            in3 => \N__11104\,
            lcout => \buart.Z_tx.bitcountZ0Z_2\,
            ltout => OPEN,
            carryin => \buart.Z_tx.un1_bitcount_cry_1\,
            carryout => \buart.Z_tx.un1_bitcount_cry_2\,
            clk => \N__29468\,
            ce => 'H',
            sr => \N__26079\
        );

    \buart.Z_tx.bitcount_3_LC_1_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101111101110"
        )
    port map (
            in0 => \N__12826\,
            in1 => \N__11092\,
            in2 => \_gnd_net_\,
            in3 => \N__11101\,
            lcout => \buart.Z_tx.bitcountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29468\,
            ce => 'H',
            sr => \N__26079\
        );

    \buart.Z_tx.bitcount_RNIVE1P1_3_LC_1_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__11518\,
            in1 => \_gnd_net_\,
            in2 => \N__11563\,
            in3 => \_gnd_net_\,
            lcout => \buart.Z_tx.bitcount_RNIVE1P1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_data_rdy_LC_1_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100000001000"
        )
    port map (
            in0 => \N__13468\,
            in1 => \N__13425\,
            in2 => \N__26158\,
            in3 => \N__12799\,
            lcout => vbuf_tx_data_rdy,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29459\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNO_0_3_LC_1_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__11519\,
            in1 => \_gnd_net_\,
            in2 => \N__11564\,
            in3 => \N__11064\,
            lcout => \buart.Z_tx.un1_bitcount_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.un1_bitcount_cry_0_0_c_RNO_LC_1_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11550\,
            in2 => \_gnd_net_\,
            in3 => \N__11517\,
            lcout => \buart.Z_tx.un1_bitcount_cry_0_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNIQOQA1_3_LC_1_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__11481\,
            in1 => \N__11076\,
            in2 => \N__11065\,
            in3 => \N__11046\,
            lcout => \buart.Z_tx.uart_busy_0_i\,
            ltout => \buart.Z_tx.uart_busy_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNI22V22_3_LC_1_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12798\,
            in2 => \N__11035\,
            in3 => \N__11516\,
            lcout => \buart.Z_tx.un1_uart_wr_i_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11120\,
            in2 => \N__11140\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_6_0_\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_2_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11152\,
            in2 => \_gnd_net_\,
            in3 => \N__11032\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_1\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_2\,
            clk => \N__29453\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_3_LC_1_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__11524\,
            in1 => \N__11161\,
            in2 => \_gnd_net_\,
            in3 => \N__11212\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_2\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_3\,
            clk => \N__29453\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_4_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11188\,
            in3 => \N__11209\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_3\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_4\,
            clk => \N__29453\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_5_LC_1_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__11525\,
            in1 => \_gnd_net_\,
            in2 => \N__11200\,
            in3 => \N__11206\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_4\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_5\,
            clk => \N__29453\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_6_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__11175\,
            in1 => \N__11523\,
            in2 => \_gnd_net_\,
            in3 => \N__11203\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29453\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_RNII048_6_LC_1_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__11196\,
            in1 => \N__11184\,
            in2 => \N__11176\,
            in3 => \N__11160\,
            lcout => OPEN,
            ltout => \buart.Z_tx.Z_baudgen.ser_clk_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_1_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__11119\,
            in1 => \N__11151\,
            in2 => \N__11143\,
            in3 => \N__11135\,
            lcout => \buart.Z_tx.ser_clk\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_1_LC_1_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__11122\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11139\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29445\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_0_LC_1_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11121\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29445\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_0_ret_29_RNO_2_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21576\,
            in1 => \N__15472\,
            in2 => \N__17565\,
            in3 => \N__15377\,
            lcout => \Lab_UT.dictrl.N_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_0_ret_29_RNO_4_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001011100000000"
        )
    port map (
            in0 => \N__20813\,
            in1 => \N__21577\,
            in2 => \N__11236\,
            in3 => \N__21110\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_17_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_0_ret_29_RNO_1_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110000"
        )
    port map (
            in0 => \N__21111\,
            in1 => \N__15473\,
            in2 => \N__11248\,
            in3 => \N__11224\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_i_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_0_ret_29_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__17137\,
            in1 => \N__24681\,
            in2 => \N__11245\,
            in3 => \N__11242\,
            lcout => \Lab_UT_dictrl_r_Sone_init17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29422\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_RNIN0MBN_1_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011100110010"
        )
    port map (
            in0 => \N__23345\,
            in1 => \N__11218\,
            in2 => \N__17929\,
            in3 => \N__17231\,
            lcout => \Lab_UT.dictrl.N_8_2\,
            ltout => \Lab_UT.dictrl.N_8_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_0_ret_29_RNO_3_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17548\,
            in2 => \N__11227\,
            in3 => \N__21575\,
            lcout => \Lab_UT.dictrl.g0_i_a8_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_RNIGHD18_0_1_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111110000"
        )
    port map (
            in0 => \N__13863\,
            in1 => \_gnd_net_\,
            in2 => \N__13834\,
            in3 => \N__18063\,
            lcout => \Lab_UT.dictrl.N_1605_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_RNO_12_1_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__18064\,
            in1 => \N__13830\,
            in2 => \_gnd_net_\,
            in3 => \N__13862\,
            lcout => \Lab_UT.dictrl.N_1605_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_RNO_7_1_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011100110010"
        )
    port map (
            in0 => \N__23376\,
            in1 => \N__17304\,
            in2 => \N__17893\,
            in3 => \N__17258\,
            lcout => \Lab_UT.dictrl.N_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_0_ret_0_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110011101111"
        )
    port map (
            in0 => \N__17260\,
            in1 => \N__24671\,
            in2 => \N__17181\,
            in3 => \N__17303\,
            lcout => \Lab_UT.dictrl.currState_i_5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29413\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_0_ret_28_RNO_4_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23375\,
            in2 => \_gnd_net_\,
            in3 => \N__17828\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.currState_0_ret_28_RNOZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_0_ret_28_RNO_2_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110100011"
        )
    port map (
            in0 => \N__17259\,
            in1 => \N__17302\,
            in2 => \N__11299\,
            in3 => \N__24669\,
            lcout => \Lab_UT.dictrl.currState_0_ret_28_RNOZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_RNO_6_1_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011100110010"
        )
    port map (
            in0 => \N__23377\,
            in1 => \N__11296\,
            in2 => \N__17894\,
            in3 => \N__17257\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_RNO_2_1_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__11290\,
            in1 => \N__15476\,
            in2 => \N__11284\,
            in3 => \N__21112\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_i_o4_4_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_RNO_0_1_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__24670\,
            in1 => \N__17572\,
            in2 => \N__11281\,
            in3 => \N__21625\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_i_o4_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010100011"
        )
    port map (
            in0 => \N__13223\,
            in1 => \N__12277\,
            in2 => \N__11278\,
            in3 => \N__15253\,
            lcout => \Lab_UT.dictrl.nextState_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29413\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.hh_0_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11275\,
            lcout => \buart.Z_rx.hhZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29405\,
            ce => 'H',
            sr => \N__26078\
        );

    \uu0.l_count_RNI04591_10_LC_2_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__11266\,
            in1 => \N__11321\,
            in2 => \N__11347\,
            in3 => \N__11395\,
            lcout => OPEN,
            ltout => \uu0.un4_l_count_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_RNI2GS72_4_LC_2_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__12513\,
            in1 => \N__12474\,
            in2 => \N__11251\,
            in3 => \N__11360\,
            lcout => OPEN,
            ltout => \uu0.un4_l_count_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_RNI8ORT6_11_LC_2_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__11437\,
            in1 => \N__11575\,
            in2 => \N__11431\,
            in3 => \N__11782\,
            lcout => \uu0.un4_l_count_0\,
            ltout => \uu0.un4_l_count_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_11_LC_2_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000011100001000"
        )
    port map (
            in0 => \N__11723\,
            in1 => \N__11425\,
            in2 => \N__11428\,
            in3 => \N__11418\,
            lcout => \uu0.l_countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29479\,
            ce => \N__12345\,
            sr => \N__26088\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_2_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__11640\,
            in1 => \N__11323\,
            in2 => \_gnd_net_\,
            in3 => \N__11397\,
            lcout => \uu0.un143_ci_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_10_LC_2_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__11725\,
            in1 => \N__11641\,
            in2 => \N__11401\,
            in3 => \N__11326\,
            lcout => \uu0.l_countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29479\,
            ce => \N__12345\,
            sr => \N__26088\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_2_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__11639\,
            in1 => \N__11322\,
            in2 => \N__11419\,
            in3 => \N__11396\,
            lcout => \uu0.un154_ci_9\,
            ltout => \uu0.un154_ci_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_14_LC_2_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__11724\,
            in1 => \N__11344\,
            in2 => \N__11365\,
            in3 => \N__11361\,
            lcout => \uu0.l_countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29479\,
            ce => \N__12345\,
            sr => \N__26088\
        );

    \uu0.l_count_9_LC_2_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11324\,
            in2 => \N__11735\,
            in3 => \N__11638\,
            lcout => \uu0.l_countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29475\,
            ce => \N__12344\,
            sr => \N__26086\
        );

    \uu0.l_count_8_LC_2_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__11325\,
            in1 => \N__11716\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uu0.l_countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29475\,
            ce => \N__12344\,
            sr => \N__26086\
        );

    \uu0.l_count_17_LC_2_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__11683\,
            in1 => \N__11604\,
            in2 => \N__11734\,
            in3 => \N__11662\,
            lcout => \uu0.l_countZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29475\,
            ce => \N__12344\,
            sr => \N__26086\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_2_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12400\,
            in1 => \N__12379\,
            in2 => \N__12433\,
            in3 => \N__11616\,
            lcout => \uu0.un110_ci\,
            ltout => \uu0.un110_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_2_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__11682\,
            in1 => \N__11603\,
            in2 => \N__11665\,
            in3 => \N__11661\,
            lcout => OPEN,
            ltout => \uu0.un220_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_18_LC_2_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11815\,
            in2 => \N__11644\,
            in3 => \N__12985\,
            lcout => \uu0.l_countZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29475\,
            ce => \N__12344\,
            sr => \N__26086\
        );

    \uu0.l_count_7_LC_2_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001010001010000"
        )
    port map (
            in0 => \N__12986\,
            in1 => \N__12493\,
            in2 => \N__11620\,
            in3 => \N__12401\,
            lcout => \uu0.l_countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29475\,
            ce => \N__12344\,
            sr => \N__26086\
        );

    \uu0.l_count_RNIRLTJ1_17_LC_2_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__11637\,
            in1 => \N__11615\,
            in2 => \N__11605\,
            in3 => \N__11588\,
            lcout => \uu0.un4_l_count_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_0_LC_2_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000011000001010"
        )
    port map (
            in0 => \N__11480\,
            in1 => \N__11569\,
            in2 => \N__12832\,
            in3 => \N__11530\,
            lcout => \buart.Z_tx.bitcountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29469\,
            ce => 'H',
            sr => \N__26084\
        );

    \uu0.delay_line_0_LC_2_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__11869\,
            in1 => \N__12523\,
            in2 => \N__11854\,
            in3 => \N__11455\,
            lcout => \uu0.delay_lineZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29469\,
            ce => 'H',
            sr => \N__26084\
        );

    \uu0.l_precount_3_LC_2_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__11457\,
            in1 => \N__11852\,
            in2 => \N__12529\,
            in3 => \N__11872\,
            lcout => \uu0.l_precountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29469\,
            ce => 'H',
            sr => \N__26084\
        );

    \uu0.l_precount_2_LC_2_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__11871\,
            in1 => \N__12525\,
            in2 => \_gnd_net_\,
            in3 => \N__11456\,
            lcout => \uu0.l_precountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29469\,
            ce => 'H',
            sr => \N__26084\
        );

    \uu0.l_precount_1_LC_2_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__12524\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11870\,
            lcout => \uu0.l_precountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29469\,
            ce => 'H',
            sr => \N__26084\
        );

    \uu0.l_precount_RNI85Q91_3_LC_2_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__11868\,
            in1 => \N__12451\,
            in2 => \N__11853\,
            in3 => \N__11830\,
            lcout => OPEN,
            ltout => \uu0.un4_l_count_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_RNI96A32_18_LC_2_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__11814\,
            in1 => \N__11803\,
            in2 => \N__11785\,
            in3 => \N__12375\,
            lcout => \uu0.un4_l_count_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_0_LC_2_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11773\,
            lcout => vbuf_tx_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__12595\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_1_LC_2_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11767\,
            lcout => vbuf_tx_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__12595\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_2_LC_2_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11761\,
            lcout => vbuf_tx_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__12595\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_3_LC_2_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11755\,
            lcout => vbuf_tx_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__12595\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_4_LC_2_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11749\,
            lcout => vbuf_tx_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__12595\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_5_LC_2_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__11743\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => vbuf_tx_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__12595\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_6_LC_2_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11953\,
            lcout => vbuf_tx_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__12595\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_7_LC_2_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11947\,
            lcout => vbuf_tx_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__12595\,
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_1_LC_2_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__11941\,
            in1 => \N__11902\,
            in2 => \_gnd_net_\,
            in3 => \N__12816\,
            lcout => \buart.Z_tx.shifterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29454\,
            ce => \N__12729\,
            sr => \N__26080\
        );

    \buart.Z_tx.shifter_0_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__12812\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11935\,
            lcout => \buart.Z_tx.shifterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29454\,
            ce => \N__12729\,
            sr => \N__26080\
        );

    \buart.Z_tx.uart_tx_LC_2_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11929\,
            in2 => \_gnd_net_\,
            in3 => \N__12819\,
            lcout => o_serial_data_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29454\,
            ce => \N__12729\,
            sr => \N__26080\
        );

    \buart.Z_tx.shifter_2_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__12813\,
            in1 => \N__11890\,
            in2 => \_gnd_net_\,
            in3 => \N__11908\,
            lcout => \buart.Z_tx.shifterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29454\,
            ce => \N__12729\,
            sr => \N__26080\
        );

    \buart.Z_tx.shifter_3_LC_2_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__11878\,
            in1 => \N__12817\,
            in2 => \_gnd_net_\,
            in3 => \N__11896\,
            lcout => \buart.Z_tx.shifterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29454\,
            ce => \N__12729\,
            sr => \N__26080\
        );

    \buart.Z_tx.shifter_4_LC_2_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__12814\,
            in1 => \N__11986\,
            in2 => \_gnd_net_\,
            in3 => \N__11884\,
            lcout => \buart.Z_tx.shifterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29454\,
            ce => \N__12729\,
            sr => \N__26080\
        );

    \buart.Z_tx.shifter_5_LC_2_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__11974\,
            in1 => \N__12818\,
            in2 => \_gnd_net_\,
            in3 => \N__11992\,
            lcout => \buart.Z_tx.shifterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29454\,
            ce => \N__12729\,
            sr => \N__26080\
        );

    \buart.Z_tx.shifter_6_LC_2_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__12815\,
            in1 => \N__12844\,
            in2 => \_gnd_net_\,
            in3 => \N__11980\,
            lcout => \buart.Z_tx.shifterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29454\,
            ce => \N__12729\,
            sr => \N__26080\
        );

    \uu2.vram_rd_clk_det_0_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13466\,
            lcout => \uu2.vram_rd_clk_detZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.vram_rd_clk_det_0C_net\,
            ce => 'H',
            sr => \N__26050\
        );

    \uu2.vram_rd_clk_det_1_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12609\,
            lcout => \uu2.vram_rd_clk_detZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.vram_rd_clk_det_0C_net\,
            ce => 'H',
            sr => \N__26050\
        );

    \uu2.l_count_3_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001001100100000"
        )
    port map (
            in0 => \N__12127\,
            in1 => \N__12938\,
            in2 => \N__13048\,
            in3 => \N__12109\,
            lcout => \uu2.l_countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29438\,
            ce => 'H',
            sr => \N__26077\
        );

    \uu2.l_count_2_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13044\,
            in2 => \_gnd_net_\,
            in3 => \N__12126\,
            lcout => \uu2.l_countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29438\,
            ce => 'H',
            sr => \N__26077\
        );

    \uu2.l_count_RNIFGGK1_3_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__12005\,
            in1 => \N__12056\,
            in2 => \N__12079\,
            in3 => \N__12107\,
            lcout => \uu2.un1_l_count_1_3\,
            ltout => \uu2.un1_l_count_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_RNI9S834_0_1_LC_2_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__13116\,
            in1 => \N__12124\,
            in2 => \N__11968\,
            in3 => \N__12091\,
            lcout => \uu2.un1_l_count_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_RNI9S834_1_LC_2_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12125\,
            in1 => \N__12145\,
            in2 => \N__11965\,
            in3 => \N__13117\,
            lcout => \uu2.un1_l_count_2_0\,
            ltout => \uu2.un1_l_count_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_4_LC_2_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000001100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12025\,
            in2 => \N__11956\,
            in3 => \N__12182\,
            lcout => \uu2.l_countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29438\,
            ce => 'H',
            sr => \N__26077\
        );

    \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12123\,
            in1 => \N__12108\,
            in2 => \N__13090\,
            in3 => \N__13115\,
            lcout => \uu2.un306_ci\,
            ltout => \uu2.un306_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_5_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101101010101010"
        )
    port map (
            in0 => \N__12057\,
            in1 => \_gnd_net_\,
            in2 => \N__12097\,
            in3 => \N__12183\,
            lcout => \uu2.l_countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29438\,
            ce => 'H',
            sr => \N__26077\
        );

    \uu2.vbuf_count.counter_gen_label_8__un350_ci_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12200\,
            in1 => \N__12006\,
            in2 => \N__12042\,
            in3 => \N__12022\,
            lcout => \uu2.un350_ci\,
            ltout => \uu2.un350_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_9_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__12078\,
            in1 => \N__12159\,
            in2 => \N__12094\,
            in3 => \N__12939\,
            lcout => \uu2.l_countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29431\,
            ce => 'H',
            sr => \N__26076\
        );

    \uu2.l_count_RNIBCGK1_0_9_LC_2_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__12198\,
            in1 => \N__12177\,
            in2 => \N__12160\,
            in3 => \N__13088\,
            lcout => \uu2.un1_l_count_1_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_8_LC_2_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12077\,
            in2 => \_gnd_net_\,
            in3 => \N__12085\,
            lcout => \uu2.l_countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29431\,
            ce => 'H',
            sr => \N__26076\
        );

    \uu2.l_count_6_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101101010101010"
        )
    port map (
            in0 => \N__12201\,
            in1 => \_gnd_net_\,
            in2 => \N__12043\,
            in3 => \N__12023\,
            lcout => \uu2.l_countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29431\,
            ce => 'H',
            sr => \N__26076\
        );

    \uu2.vbuf_count.counter_gen_label_6__un328_ci_3_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__12181\,
            in1 => \N__12058\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uu2.vbuf_count.un328_ci_3\,
            ltout => \uu2.vbuf_count.un328_ci_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_7_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__12202\,
            in1 => \N__12007\,
            in2 => \N__12028\,
            in3 => \N__12024\,
            lcout => \uu2.l_countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29431\,
            ce => 'H',
            sr => \N__26076\
        );

    \uu2.l_count_RNIBCGK1_9_LC_2_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__13089\,
            in1 => \N__12199\,
            in2 => \N__12184\,
            in3 => \N__12158\,
            lcout => \uu2.un1_l_count_2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_0_rep2_RNIOBFP3_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__24878\,
            in1 => \N__27790\,
            in2 => \N__20950\,
            in3 => \N__27542\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_8_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_RNIA5707_2_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011001000"
        )
    port map (
            in0 => \N__25020\,
            in1 => \N__12214\,
            in2 => \N__12139\,
            in3 => \N__12133\,
            lcout => \Lab_UT.dictrl.N_23_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__g0_13_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__20949\,
            in1 => \N__27789\,
            in2 => \_gnd_net_\,
            in3 => \N__27541\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_20_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__g0_5_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011111001111"
        )
    port map (
            in0 => \N__21245\,
            in1 => \N__23826\,
            in2 => \N__12136\,
            in3 => \N__17112\,
            lcout => \Lab_UT.dictrl.N_30_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_RNIKTU5_2_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15541\,
            in2 => \_gnd_net_\,
            in3 => \N__23326\,
            lcout => \Lab_UT.dictrl.G_19_0_a7_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_0_ret_21_RNI40BJ2_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__27296\,
            in1 => \N__20361\,
            in2 => \_gnd_net_\,
            in3 => \N__24005\,
            lcout => \Lab_UT.dictrl.N_9_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_3_3_rep1_RNIO9JG3_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__20360\,
            in1 => \N__27297\,
            in2 => \N__14269\,
            in3 => \N__23327\,
            lcout => \Lab_UT.dictrl.G_30_0_a7_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_fast_RNI13TV_0_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__25019\,
            in1 => \N__17861\,
            in2 => \N__24897\,
            in3 => \N__14500\,
            lcout => \Lab_UT.dictrl.G_30_0_a7_4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_0_ret_29_RNIK6A94_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__27561\,
            in1 => \N__27809\,
            in2 => \N__12253\,
            in3 => \N__23341\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_31_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_0_ret_29_RNINPDOC_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110010"
        )
    port map (
            in0 => \N__12244\,
            in1 => \N__12271\,
            in2 => \N__12238\,
            in3 => \N__12220\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.G_30_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_0_ret_21_RNI66NNS_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__12265\,
            in1 => \N__12235\,
            in2 => \N__12229\,
            in3 => \N__21133\,
            lcout => \Lab_UT.dictrl.nextStateZ0Z_1\,
            ltout => \Lab_UT.dictrl.nextStateZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_0_ret_21_RNIAVHPS_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12226\,
            in3 => \N__24680\,
            lcout => \Lab_UT.dictrl.N_10ctr\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_3_3_rep1_RNIPTVF_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17860\,
            in2 => \_gnd_net_\,
            in3 => \N__20334\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.G_30_0_a7_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_RNIO37J1_1_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010001000"
        )
    port map (
            in0 => \N__23343\,
            in1 => \N__13216\,
            in2 => \N__12223\,
            in3 => \N__14268\,
            lcout => \Lab_UT.dictrl.G_30_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_RNI1O2A_1_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17859\,
            in2 => \_gnd_net_\,
            in3 => \N__23340\,
            lcout => \Lab_UT.dictrl.G_30_0_a7_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_RNI0P25D_1_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000011110100"
        )
    port map (
            in0 => \N__23342\,
            in1 => \N__17862\,
            in2 => \N__15157\,
            in3 => \N__12208\,
            lcout => \Lab_UT.dictrl.currState_2_RNI0P25DZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__g0_0_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010001000"
        )
    port map (
            in0 => \N__25045\,
            in1 => \N__13864\,
            in2 => \N__24899\,
            in3 => \N__15336\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.i8_mux_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__g0_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__17888\,
            in1 => \_gnd_net_\,
            in2 => \N__12280\,
            in3 => \N__17261\,
            lcout => \Lab_UT.dictrl.i7_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_RNIJ59B3_2_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__25041\,
            in1 => \N__17886\,
            in2 => \N__24898\,
            in3 => \N__27543\,
            lcout => \Lab_UT.dictrl.N_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_1_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24673\,
            in2 => \_gnd_net_\,
            in3 => \N__20622\,
            lcout => \Lab_UT_dictrl_currState_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29406\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_ret_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111010111111"
        )
    port map (
            in0 => \N__24672\,
            in1 => \N__18061\,
            in2 => \N__15583\,
            in3 => \N__14025\,
            lcout => \Lab_UT.dictrl.currState_i_5_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29406\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_fast_0_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24674\,
            in2 => \_gnd_net_\,
            in3 => \N__21109\,
            lcout => \Lab_UT.dictrl.currState_fast_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29406\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_RNITUPT_2_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__23344\,
            in1 => \N__23814\,
            in2 => \N__25048\,
            in3 => \N__17887\,
            lcout => \Lab_UT.dictrl.G_30_0_a7_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_3_3_rep1_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__21608\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24675\,
            lcout => \Lab_UT.dictrl.currState_3_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29406\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_0_ret_21_RNIUL8L_0_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__23825\,
            in1 => \N__18060\,
            in2 => \_gnd_net_\,
            in3 => \N__24007\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_11_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_RNIKSEU7_0_0_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__21234\,
            in1 => \N__12313\,
            in2 => \N__12256\,
            in3 => \N__27787\,
            lcout => \Lab_UT.dictrl.N_5_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_0_ret_24_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__17567\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15483\,
            lcout => \Lab_UT.dictrl.r_dicLdMtens22_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29399\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_RNIHF8J71_1_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010000000"
        )
    port map (
            in0 => \N__12325\,
            in1 => \N__21607\,
            in2 => \N__17892\,
            in3 => \N__17262\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_RNIDEJTG4_1_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__17566\,
            in1 => \N__15482\,
            in2 => \N__12319\,
            in3 => \N__21098\,
            lcout => \Lab_UT.dictrl.N_7_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_3_RNIR9C03_3_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__18058\,
            in1 => \N__23824\,
            in2 => \_gnd_net_\,
            in3 => \N__27298\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_8_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_ret_5_RNIN6436_0_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011110000"
        )
    port map (
            in0 => \N__24888\,
            in1 => \N__18059\,
            in2 => \N__12316\,
            in3 => \N__27552\,
            lcout => \Lab_UT.dictrl.N_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_ret_RNI7FNU_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010101010"
        )
    port map (
            in0 => \N__12307\,
            in1 => \N__23860\,
            in2 => \_gnd_net_\,
            in3 => \N__24889\,
            lcout => \Lab_UT.dictrl.currState_ret_RNI7FNUZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_fast_RNIT3362_0_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14501\,
            in1 => \N__17428\,
            in2 => \N__24901\,
            in3 => \N__12535\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.G_19_0_a7_4_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_fast_RNIOKOT3_0_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12541\,
            in1 => \N__18187\,
            in2 => \N__12301\,
            in3 => \N__17668\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_0_rep2_RNI0FS1A_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110010"
        )
    port map (
            in0 => \N__12547\,
            in1 => \N__24477\,
            in2 => \N__12298\,
            in3 => \N__12286\,
            lcout => \Lab_UT.dictrl.G_19_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_ret_5_RNIIF461_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__18057\,
            in1 => \N__17855\,
            in2 => \N__24900\,
            in3 => \N__12295\,
            lcout => \Lab_UT.dictrl.G_19_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_0_rep2_RNI5U4U_LC_2_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18056\,
            in1 => \N__17854\,
            in2 => \N__20940\,
            in3 => \N__20369\,
            lcout => \Lab_UT.dictrl.G_19_0_a7_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_6_rep1_RNI4H7E_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__23422\,
            in1 => \N__22000\,
            in2 => \N__17910\,
            in3 => \N__21415\,
            lcout => \G_19_0_a7_4_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_4_rep1_RNI7DDT_LC_2_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21841\,
            in2 => \_gnd_net_\,
            in3 => \N__21444\,
            lcout => \G_19_0_a7_4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.hh_1_LC_2_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14292\,
            lcout => \buart.Z_rx.hhZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29383\,
            ce => 'H',
            sr => \N__26087\
        );

    \uu0.l_precount_0_LC_4_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12512\,
            lcout => \uu0.l_precountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29470\,
            ce => 'H',
            sr => \N__26093\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_4_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12426\,
            in2 => \_gnd_net_\,
            in3 => \N__12373\,
            lcout => \uu0.un99_ci_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_5_LC_4_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__12411\,
            in1 => \N__12481\,
            in2 => \_gnd_net_\,
            in3 => \N__12450\,
            lcout => \uu0.l_countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29455\,
            ce => \N__12346\,
            sr => \N__26089\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_4_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12480\,
            in2 => \_gnd_net_\,
            in3 => \N__12449\,
            lcout => \uu0.un88_ci_3\,
            ltout => \uu0.un88_ci_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_6_LC_4_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__12374\,
            in1 => \N__12412\,
            in2 => \N__12382\,
            in3 => \N__13007\,
            lcout => \uu0.l_countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29455\,
            ce => \N__12346\,
            sr => \N__26089\
        );

    \uu2.mem0.ram512X8_inst_RNO_7_LC_4_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__16645\,
            in1 => \N__16177\,
            in2 => \_gnd_net_\,
            in3 => \N__18775\,
            lcout => \uu2.mem0.w_addr_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vram_rd_clk_det_RNI95711_1_LC_4_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__12625\,
            in1 => \N__12613\,
            in2 => \_gnd_net_\,
            in3 => \N__26144\,
            lcout => \uu2.vram_rd_clk_det_RNI95711Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Mones_subtractor.q20_0_i_LC_4_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__26145\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26929\,
            lcout => \Lab_UT.didp.q20_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.uu0.l_count_RNIP43E_13_LC_4_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16033\,
            in2 => \_gnd_net_\,
            in3 => \N__16009\,
            lcout => \Lab_UT.uu0.un4_l_count_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_12_LC_4_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__12666\,
            in1 => \N__22639\,
            in2 => \_gnd_net_\,
            in3 => \N__18798\,
            lcout => \uu2.mem0.w_data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_13_LC_4_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__18799\,
            in1 => \N__12568\,
            in2 => \_gnd_net_\,
            in3 => \N__22618\,
            lcout => \uu2.mem0.w_data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIOA9K6_8_LC_4_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000100"
        )
    port map (
            in0 => \N__16399\,
            in1 => \N__13024\,
            in2 => \N__16057\,
            in3 => \N__18864\,
            lcout => \uu2.N_37\,
            ltout => \uu2.N_37_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_11_LC_4_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111011000"
        )
    port map (
            in0 => \N__18801\,
            in1 => \N__22834\,
            in2 => \N__12562\,
            in3 => \N__12870\,
            lcout => \uu2.mem0.w_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_9_LC_4_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111010"
        )
    port map (
            in0 => \N__12667\,
            in1 => \N__22666\,
            in2 => \N__12874\,
            in3 => \N__18802\,
            lcout => \uu2.mem0.w_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI7QIF3_8_LC_4_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__13023\,
            in1 => \N__16053\,
            in2 => \_gnd_net_\,
            in3 => \N__16398\,
            lcout => OPEN,
            ltout => \uu2.N_51_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIEK5V6_0_LC_4_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18865\,
            in2 => \N__12670\,
            in3 => \N__19494\,
            lcout => \uu2.N_34\,
            ltout => \uu2.N_34_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_8_LC_4_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__18800\,
            in1 => \_gnd_net_\,
            in2 => \N__12658\,
            in3 => \N__25682\,
            lcout => \uu2.mem0.w_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIASLS1_4_LC_4_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110010101101010"
        )
    port map (
            in0 => \N__14919\,
            in1 => \N__16512\,
            in2 => \N__14590\,
            in3 => \N__16275\,
            lcout => OPEN,
            ltout => \uu2.bitmap_pmux_sn_m15_0_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIIO5V6_2_LC_4_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101010100000"
        )
    port map (
            in0 => \N__12862\,
            in1 => \N__12646\,
            in2 => \N__12649\,
            in3 => \N__14589\,
            lcout => \uu2.bitmap_pmux_sn_i7_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIV2MM2_2_LC_4_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000010000"
        )
    port map (
            in0 => \N__14918\,
            in1 => \N__19493\,
            in2 => \N__13525\,
            in3 => \N__16274\,
            lcout => \uu2.bitmap_pmux_sn_N_65\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI03P31_4_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011000110011"
        )
    port map (
            in0 => \N__16513\,
            in1 => \N__14920\,
            in2 => \_gnd_net_\,
            in3 => \N__16129\,
            lcout => OPEN,
            ltout => \uu2.bitmap_pmux_sn_m24_0_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIEFIL2_0_LC_4_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001100000000110"
        )
    port map (
            in0 => \N__14585\,
            in1 => \N__19492\,
            in2 => \N__12640\,
            in3 => \N__16273\,
            lcout => OPEN,
            ltout => \uu2.bitmap_pmux_sn_i5_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI0HFE3_8_LC_4_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16787\,
            in2 => \N__12637\,
            in3 => \N__16643\,
            lcout => OPEN,
            ltout => \uu2.bitmap_pmux_29_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI649331_8_LC_4_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001000000"
        )
    port map (
            in0 => \N__12883\,
            in1 => \N__13705\,
            in2 => \N__12877\,
            in3 => \N__13501\,
            lcout => \uu2.bitmap_pmux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI12TI1_5_LC_4_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000010100000"
        )
    port map (
            in0 => \N__16549\,
            in1 => \N__16786\,
            in2 => \N__16447\,
            in3 => \N__16642\,
            lcout => \uu2.bitmap_pmux_sn_N_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_7_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12830\,
            in2 => \N__12745\,
            in3 => \N__12856\,
            lcout => \buart.Z_tx.shifterZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29432\,
            ce => \N__12736\,
            sr => \N__26082\
        );

    \buart.Z_tx.shifter_8_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__12831\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12757\,
            lcout => \buart.Z_tx.shifterZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29432\,
            ce => \N__12736\,
            sr => \N__26082\
        );

    \uu0.delay_line_RNILLLG7_1_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__12892\,
            in1 => \N__12915\,
            in2 => \_gnd_net_\,
            in3 => \N__13011\,
            lcout => \uu0.un11_l_count_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNIUEOT_58_LC_4_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__16816\,
            in1 => \N__19084\,
            in2 => \_gnd_net_\,
            in3 => \N__16788\,
            lcout => \uu2.N_161\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_6_LC_4_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__16789\,
            in1 => \N__16159\,
            in2 => \_gnd_net_\,
            in3 => \N__18786\,
            lcout => \uu2.mem0.w_addr_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_0_LC_4_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__16132\,
            in1 => \N__18973\,
            in2 => \_gnd_net_\,
            in3 => \N__18785\,
            lcout => \uu2.mem0.w_addr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_nesr_RNI4JSO_1_LC_4_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19487\,
            in2 => \_gnd_net_\,
            in3 => \N__16130\,
            lcout => \uu2.N_31_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI25P31_8_LC_4_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__16131\,
            in1 => \_gnd_net_\,
            in2 => \N__19498\,
            in3 => \N__16644\,
            lcout => \uu2.w_data_displaying_2_i_a2_i_a3_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.sec_clk_LC_4_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26794\,
            in2 => \_gnd_net_\,
            in3 => \N__13012\,
            lcout => \o_One_Sec_Pulse\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29423\,
            ce => 'H',
            sr => \N__26081\
        );

    \uu2.l_count_1_LC_4_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13078\,
            in2 => \_gnd_net_\,
            in3 => \N__13114\,
            lcout => \uu2.l_countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29423\,
            ce => 'H',
            sr => \N__26081\
        );

    \uu2.l_count_0_LC_4_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__13079\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uu2.l_countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29423\,
            ce => 'H',
            sr => \N__26081\
        );

    \uu2.vram_rd_clk_LC_4_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13450\,
            in2 => \_gnd_net_\,
            in3 => \N__12940\,
            lcout => \uu2.vram_rd_clkZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29423\,
            ce => 'H',
            sr => \N__26081\
        );

    \Lab_UT.uu0.delay_line_1_LC_4_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22153\,
            lcout => \Lab_UT.uu0.delay_lineZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29423\,
            ce => 'H',
            sr => \N__26081\
        );

    \uu0.delay_line_1_LC_4_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12919\,
            lcout => \uu0.delay_lineZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29423\,
            ce => 'H',
            sr => \N__26081\
        );

    \Lab_UT.dictrl.currState_ret_2_LC_4_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__24626\,
            in1 => \N__20814\,
            in2 => \_gnd_net_\,
            in3 => \N__21624\,
            lcout => \Lab_UT.dictrl.r_dicLdMtens23_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29414\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_0_LC_4_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24627\,
            in2 => \_gnd_net_\,
            in3 => \N__21108\,
            lcout => \Lab_UT.dictrl.currStateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29414\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.sec_clkD_RNISDHD_LC_4_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__26784\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26748\,
            lcout => \oneSecStrb\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.sec_clkD_LC_4_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26785\,
            lcout => \uu0_sec_clkD\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29414\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_count.counter_gen_label_2__un284_ci_LC_4_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13113\,
            in2 => \_gnd_net_\,
            in3 => \N__13077\,
            lcout => \uu2.un284_ci\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_ness_RNO_0_6_LC_4_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16465\,
            in2 => \_gnd_net_\,
            in3 => \N__16375\,
            lcout => \uu2.N_48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.rst_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19191\,
            lcout => rst,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29407\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_ret_RNI5RB74_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__27295\,
            in1 => \N__13896\,
            in2 => \_gnd_net_\,
            in3 => \N__27792\,
            lcout => \Lab_UT.dictrl.dicLdAMtens_rst\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__m8_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__20392\,
            in1 => \N__14179\,
            in2 => \_gnd_net_\,
            in3 => \N__14161\,
            lcout => \Lab_UT.dictrl.N_9\,
            ltout => \Lab_UT.dictrl.N_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_RNINHPTJ_1_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000010100010"
        )
    port map (
            in0 => \N__13948\,
            in1 => \N__17916\,
            in2 => \N__13030\,
            in3 => \N__20284\,
            lcout => \Lab_UT.dictrl.N_19_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_RNIR9C03_2_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__25008\,
            in1 => \N__23430\,
            in2 => \N__23833\,
            in3 => \N__27294\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_21_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_ret_5_RNIN6436_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011110000"
        )
    port map (
            in0 => \N__24864\,
            in1 => \N__18014\,
            in2 => \N__13027\,
            in3 => \N__27551\,
            lcout => \Lab_UT.dictrl.N_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__g0_0_0_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14101\,
            in2 => \_gnd_net_\,
            in3 => \N__27293\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__g0_1_LC_4_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100010001000"
        )
    port map (
            in0 => \N__23972\,
            in1 => \N__23827\,
            in2 => \N__13138\,
            in3 => \N__27791\,
            lcout => \Lab_UT.dictrl.N_23_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__m21_mb_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__13144\,
            in1 => \N__23818\,
            in2 => \N__25039\,
            in3 => \N__14455\,
            lcout => \Lab_UT.dictrl.i8_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_0_ret_21_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__13192\,
            in1 => \N__13183\,
            in2 => \N__13126\,
            in3 => \N__13168\,
            lcout => \Lab_UT.dictrl.currState_i_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29400\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_0_ret_1_RNINTRN4_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__27747\,
            in1 => \N__23898\,
            in2 => \_gnd_net_\,
            in3 => \N__27277\,
            lcout => \Lab_UT.dictrl.dicLdAStens_rst\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_RNIA8EV3_0_1_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011110101"
        )
    port map (
            in0 => \N__23381\,
            in1 => \N__13252\,
            in2 => \N__13237\,
            in3 => \N__27745\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_1611_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_RNIFHD18_1_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18006\,
            in2 => \N__13135\,
            in3 => \N__13132\,
            lcout => \Lab_UT.dictrl.N_1605_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_3_RNI3HN91_3_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__14209\,
            in1 => \N__23817\,
            in2 => \_gnd_net_\,
            in3 => \N__18115\,
            lcout => \Lab_UT.dictrl.G_28_0_a5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_RNI0LLB7_0_LC_4_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__27746\,
            in1 => \N__15349\,
            in2 => \N__21244\,
            in3 => \N__27276\,
            lcout => \Lab_UT.dictrl.N_8_3\,
            ltout => \Lab_UT.dictrl.N_8_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_RNIQ7IPD1_0_LC_4_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__13191\,
            in1 => \N__13182\,
            in2 => \N__13174\,
            in3 => \N__13167\,
            lcout => \Lab_UT.dictrl.N_6ctr\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_0_rep2_RNIBGCI9_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__13153\,
            in1 => \N__14107\,
            in2 => \N__13279\,
            in3 => \N__13159\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.currState_2_0_rep2_RNIBGCIZ0Z9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_RNI0GB6H_0_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000011000100"
        )
    port map (
            in0 => \N__18111\,
            in1 => \N__14205\,
            in2 => \N__13171\,
            in3 => \N__13981\,
            lcout => \Lab_UT.dictrl.G_28_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_0_rep2_RNIKH8P2_LC_4_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100110011"
        )
    port map (
            in0 => \N__20936\,
            in1 => \N__29073\,
            in2 => \_gnd_net_\,
            in3 => \N__27248\,
            lcout => \Lab_UT.dictrl.currState_2_0_rep2_RNIKH8PZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_RNI0KKK6_0_LC_4_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001110010"
        )
    port map (
            in0 => \N__18041\,
            in1 => \N__24813\,
            in2 => \N__14008\,
            in3 => \N__13243\,
            lcout => \Lab_UT.dictrl.N_1609_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_RNIS6CF1_5_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__28981\,
            in1 => \N__24448\,
            in2 => \_gnd_net_\,
            in3 => \N__27731\,
            lcout => \shifter_RNIS6CF1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__g0_4_LC_4_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010110011101100"
        )
    port map (
            in0 => \N__27247\,
            in1 => \N__20937\,
            in2 => \N__27788\,
            in3 => \N__27517\,
            lcout => \Lab_UT.dictrl.N_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__m21_rn_1_0_LC_4_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__20935\,
            in1 => \N__27730\,
            in2 => \_gnd_net_\,
            in3 => \N__27249\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.m21_rn_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__m21_rn_LC_4_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001011111010"
        )
    port map (
            in0 => \N__25012\,
            in1 => \N__24814\,
            in2 => \N__13147\,
            in3 => \N__15320\,
            lcout => \Lab_UT.dictrl.m21_rn_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_ret_5_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0001101110111011"
        )
    port map (
            in0 => \N__18046\,
            in1 => \N__13957\,
            in2 => \N__13974\,
            in3 => \N__17915\,
            lcout => \Lab_UT.dictrl.currState_i_5_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29389\,
            ce => 'H',
            sr => \N__26064\
        );

    \Lab_UT.dictrl.currState_2_0_rep1_RNI3BNS2_LC_4_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__27483\,
            in1 => \N__24802\,
            in2 => \_gnd_net_\,
            in3 => \N__14088\,
            lcout => \Lab_UT.dictrl.g1_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__g0_17_LC_4_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110011111100"
        )
    port map (
            in0 => \N__27645\,
            in1 => \N__14347\,
            in2 => \N__14096\,
            in3 => \N__27212\,
            lcout => \Lab_UT.dictrl.N_13_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__g0_18_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111011001100"
        )
    port map (
            in0 => \N__27210\,
            in1 => \N__14087\,
            in2 => \N__27510\,
            in3 => \N__27646\,
            lcout => \Lab_UT.dictrl.N_7_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__m4_LC_4_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101100011111000"
        )
    port map (
            in0 => \N__27643\,
            in1 => \N__27475\,
            in2 => \N__14095\,
            in3 => \N__27209\,
            lcout => \Lab_UT.dictrl.N_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__m6_LC_4_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111011001100"
        )
    port map (
            in0 => \N__27211\,
            in1 => \N__14083\,
            in2 => \N__27511\,
            in3 => \N__27644\,
            lcout => \Lab_UT.dictrl.N_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__m19_LC_4_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000010000000"
        )
    port map (
            in0 => \N__27647\,
            in1 => \N__27482\,
            in2 => \N__14097\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.dictrl.N_20\,
            ltout => \Lab_UT.dictrl.N_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_RNIA8EV3_1_LC_4_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000111111"
        )
    port map (
            in0 => \N__13233\,
            in1 => \N__24803\,
            in2 => \N__13195\,
            in3 => \N__23431\,
            lcout => \Lab_UT.dictrl.nextState_RNIA8EV3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.decoder.de_littleA_2_0_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21389\,
            in1 => \N__21441\,
            in2 => \N__21767\,
            in3 => \N__21683\,
            lcout => \Lab_UT.dictrl.decoder.de_littleA_2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.decoder.de_num_0_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000101010"
        )
    port map (
            in0 => \N__14223\,
            in1 => \N__21749\,
            in2 => \N__21698\,
            in3 => \N__21392\,
            lcout => \Lab_UT.dictrl.de_num_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.decoder.de_num0to5_1_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100000000"
        )
    port map (
            in0 => \N__21391\,
            in1 => \N__21685\,
            in2 => \N__21766\,
            in3 => \N__14222\,
            lcout => \Lab_UT.dictrl.de_num0to5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.decoder.g0_1_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21390\,
            in2 => \_gnd_net_\,
            in3 => \N__21352\,
            lcout => \Lab_UT.dictrl.decoder.g0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.decoder.g0_5_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21756\,
            in1 => \N__21684\,
            in2 => \N__21999\,
            in3 => \N__21936\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.decoder.g0Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.decoder.g0_6_LC_4_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__25372\,
            in1 => \N__25272\,
            in2 => \N__13264\,
            in3 => \N__13261\,
            lcout => \Lab_UT.dictrl.g0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__g0_21_LC_4_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__21222\,
            in1 => \N__27773\,
            in2 => \N__18400\,
            in3 => \N__27246\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_36_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__g0_20_LC_4_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__14239\,
            in1 => \N__15304\,
            in2 => \N__13255\,
            in3 => \N__23815\,
            lcout => \Lab_UT.dictrl.N_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_4_rep1_LC_4_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24415\,
            lcout => bu_rx_data_4_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29380\,
            ce => \N__25428\,
            sr => \N__26090\
        );

    \buart.Z_rx.shifter_1_rep1_LC_4_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28596\,
            lcout => bu_rx_data_1_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29380\,
            ce => \N__25428\,
            sr => \N__26090\
        );

    \buart.Z_rx.shifter_3_rep1_LC_4_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25279\,
            lcout => bu_rx_data_3_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29380\,
            ce => \N__25428\,
            sr => \N__26090\
        );

    \buart.Z_rx.shifter_fast_7_LC_4_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__21877\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_fast_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29380\,
            ce => \N__25428\,
            sr => \N__26090\
        );

    \buart.Z_rx.shifter_4_LC_4_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__24416\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29380\,
            ce => \N__25428\,
            sr => \N__26090\
        );

    \buart.Z_rx.shifter_2_rep1_LC_4_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__28982\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_2_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29380\,
            ce => \N__25428\,
            sr => \N__26090\
        );

    \Lab_UT.dictrl.nextState_1_3_0__m7_LC_4_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011111100"
        )
    port map (
            in0 => \N__27716\,
            in1 => \N__24004\,
            in2 => \N__14437\,
            in3 => \N__14224\,
            lcout => \Lab_UT.dictrl.N_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_3_3_rep1_RNIM4AP_LC_4_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__25344\,
            in1 => \N__28613\,
            in2 => \_gnd_net_\,
            in3 => \N__20370\,
            lcout => OPEN,
            ltout => \G_28_0_a5_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_RNI1D8L1_4_LC_4_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__28817\,
            in1 => \N__24266\,
            in2 => \N__13282\,
            in3 => \N__25273\,
            lcout => \shifter_RNI1D8L1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_6_LC_4_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__25345\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29375\,
            ce => \N__25425\,
            sr => \N__26092\
        );

    \buart.Z_rx.shifter_fast_6_LC_4_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__25346\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_fast_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29375\,
            ce => \N__25425\,
            sr => \N__26092\
        );

    \buart.Z_rx.shifter_7_LC_4_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21871\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29375\,
            ce => \N__25425\,
            sr => \N__26092\
        );

    \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_4_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14415\,
            in2 => \N__13297\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_16_0_\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_4_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13308\,
            in2 => \_gnd_net_\,
            in3 => \N__13267\,
            lcout => \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.Z_baudgen.un5_counter_cry_1\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_3_LC_4_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__15926\,
            in1 => \N__14428\,
            in2 => \_gnd_net_\,
            in3 => \N__13339\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \buart.Z_rx.Z_baudgen.un5_counter_cry_2\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_3\,
            clk => \N__29373\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_4_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14380\,
            in3 => \N__13336\,
            lcout => \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.Z_baudgen.un5_counter_cry_3\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_5_LC_4_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000100"
        )
    port map (
            in0 => \N__15925\,
            in1 => \N__13329\,
            in2 => \N__15625\,
            in3 => \N__13333\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29373\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_RNI4IE3_5_LC_4_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__14375\,
            in1 => \N__13307\,
            in2 => \N__13330\,
            in3 => \N__13292\,
            lcout => \buart.Z_rx.Z_baudgen.ser_clk_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_2_LC_4_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__13309\,
            in1 => \N__15924\,
            in2 => \N__13318\,
            in3 => \N__15624\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29373\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_1_LC_4_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__15923\,
            in1 => \N__14416\,
            in2 => \_gnd_net_\,
            in3 => \N__13296\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29373\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_addr_2_LC_5_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__13626\,
            in1 => \N__13589\,
            in2 => \N__13662\,
            in3 => \N__25133\,
            lcout => \uu2.r_addrZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29447\,
            ce => 'H',
            sr => \N__26068\
        );

    \uu2.r_addr_1_LC_5_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__25132\,
            in1 => \_gnd_net_\,
            in2 => \N__13593\,
            in3 => \N__13625\,
            lcout => \uu2.r_addrZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29447\,
            ce => 'H',
            sr => \N__26068\
        );

    \uu2.trig_rd_det_RNINBDQ_1_LC_5_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25131\,
            in2 => \_gnd_net_\,
            in3 => \N__26150\,
            lcout => \uu2.trig_rd_is_det_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.trig_rd_det_RNIJIIO_1_LC_5_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13474\,
            in2 => \_gnd_net_\,
            in3 => \N__13407\,
            lcout => \uu2.trig_rd_is_det\,
            ltout => \uu2.trig_rd_is_det_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_addr_0_LC_5_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13477\,
            in3 => \N__13585\,
            lcout => \uu2.r_addrZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29447\,
            ce => 'H',
            sr => \N__26068\
        );

    \uu2.trig_rd_det_1_LC_5_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13408\,
            lcout => \uu2.trig_rd_detZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29447\,
            ce => 'H',
            sr => \N__26068\
        );

    \uu2.trig_rd_det_0_LC_5_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13467\,
            in2 => \_gnd_net_\,
            in3 => \N__13426\,
            lcout => \uu2.trig_rd_detZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29447\,
            ce => 'H',
            sr => \N__26068\
        );

    \uu2.vbuf_raddr.counter_gen_label_8__un448_ci_0_LC_5_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13355\,
            in2 => \_gnd_net_\,
            in3 => \N__13684\,
            lcout => \uu2.vbuf_raddr.un448_ci_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_raddr.counter_gen_label_6__un426_ci_3_LC_5_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__22793\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25109\,
            lcout => \uu2.vbuf_raddr.un426_ci_3\,
            ltout => \uu2.vbuf_raddr.un426_ci_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_addr_esr_8_LC_5_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__13383\,
            in1 => \N__13399\,
            in2 => \N__13393\,
            in3 => \N__25160\,
            lcout => \uu2.r_addrZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29439\,
            ce => \N__13534\,
            sr => \N__26066\
        );

    \uu2.r_addr_esr_7_LC_5_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__25161\,
            in1 => \N__13356\,
            in2 => \N__13692\,
            in3 => \N__13369\,
            lcout => \uu2.r_addrZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29439\,
            ce => \N__13534\,
            sr => \N__26066\
        );

    \uu2.vbuf_raddr.counter_gen_label_4__un404_ci_LC_5_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__13654\,
            in1 => \N__13623\,
            in2 => \N__13556\,
            in3 => \N__13583\,
            lcout => \uu2.un404_ci_0\,
            ltout => \uu2.un404_ci_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_addr_esr_6_LC_5_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__13688\,
            in1 => \N__22807\,
            in2 => \N__13699\,
            in3 => \N__25110\,
            lcout => \uu2.r_addrZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29439\,
            ce => \N__13534\,
            sr => \N__26066\
        );

    \uu2.r_addr_esr_3_LC_5_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__13655\,
            in1 => \N__13624\,
            in2 => \N__13557\,
            in3 => \N__13584\,
            lcout => \uu2.r_addrZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29439\,
            ce => \N__13534\,
            sr => \N__26066\
        );

    \uu2.w_addr_displaying_RNI12TI1_0_5_LC_5_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001101001000"
        )
    port map (
            in0 => \N__16545\,
            in1 => \N__16768\,
            in2 => \N__16442\,
            in3 => \N__16627\,
            lcout => \uu2.bitmap_pmux_sn_N_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNIHNN91_40_LC_5_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110001110111"
        )
    port map (
            in0 => \N__13762\,
            in1 => \N__16257\,
            in2 => \N__13756\,
            in3 => \N__16640\,
            lcout => OPEN,
            ltout => \uu2.bitmap_pmux_26_bm_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNI1PH82_34_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111000001110"
        )
    port map (
            in0 => \N__16258\,
            in1 => \N__13483\,
            in2 => \N__13516\,
            in3 => \N__14950\,
            lcout => \uu2.bitmap_RNI1PH82Z0Z_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI2NHS5_8_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000011111101"
        )
    port map (
            in0 => \N__16259\,
            in1 => \N__16641\,
            in2 => \N__13513\,
            in3 => \N__14632\,
            lcout => OPEN,
            ltout => \uu2.N_400_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIB4NVD_4_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14626\,
            in2 => \N__13504\,
            in3 => \N__13489\,
            lcout => \uu2.N_409\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNIPUBH6_34_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__14929\,
            in1 => \N__13495\,
            in2 => \_gnd_net_\,
            in3 => \N__14608\,
            lcout => \uu2.N_404\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_290_LC_5_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101010101010"
        )
    port map (
            in0 => \N__19888\,
            in1 => \N__17056\,
            in2 => \N__15064\,
            in3 => \N__16870\,
            lcout => \uu2.bitmapZ0Z_290\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_290C_net\,
            ce => 'H',
            sr => \N__26041\
        );

    \uu2.bitmap_40_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__15118\,
            in1 => \N__19889\,
            in2 => \_gnd_net_\,
            in3 => \N__14863\,
            lcout => \uu2.bitmapZ0Z_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_290C_net\,
            ce => 'H',
            sr => \N__26041\
        );

    \uu2.bitmap_296_LC_5_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011110000"
        )
    port map (
            in0 => \N__14854\,
            in1 => \_gnd_net_\,
            in2 => \N__19897\,
            in3 => \N__15117\,
            lcout => \uu2.bitmapZ0Z_296\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_290C_net\,
            ce => 'H',
            sr => \N__26041\
        );

    \uu2.bitmap_RNIIOM81_66_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001111"
        )
    port map (
            in0 => \N__13735\,
            in1 => \N__19436\,
            in2 => \N__14980\,
            in3 => \N__16769\,
            lcout => OPEN,
            ltout => \uu2.bitmap_pmux_25_am_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNIM7D32_69_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__19437\,
            in1 => \N__13744\,
            in2 => \N__13747\,
            in3 => \N__14965\,
            lcout => \uu2.bitmap_RNIM7D32Z0Z_69\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_197_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101110"
        )
    port map (
            in0 => \N__19884\,
            in1 => \N__15060\,
            in2 => \N__17071\,
            in3 => \N__16846\,
            lcout => \uu2.bitmapZ0Z_197\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_197C_net\,
            ce => 'H',
            sr => \N__26039\
        );

    \uu2.bitmap_66_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__15059\,
            in1 => \N__19885\,
            in2 => \_gnd_net_\,
            in3 => \N__16894\,
            lcout => \uu2.bitmapZ0Z_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_197C_net\,
            ce => 'H',
            sr => \N__26039\
        );

    \uu2.bitmap_RNI2JA82_212_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110111000"
        )
    port map (
            in0 => \N__16699\,
            in1 => \N__14659\,
            in2 => \N__16669\,
            in3 => \N__16770\,
            lcout => OPEN,
            ltout => \uu2.bitmap_RNI2JA82Z0Z_212_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_nesr_RNIEE9K5_3_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101100111"
        )
    port map (
            in0 => \N__13725\,
            in1 => \N__16267\,
            in2 => \N__13729\,
            in3 => \N__13768\,
            lcout => OPEN,
            ltout => \uu2.bitmap_pmux_27_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNI9MSLA_69_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__13726\,
            in1 => \N__13714\,
            in2 => \N__13708\,
            in3 => \N__19369\,
            lcout => \uu2.N_407\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment3.segmentUQ_0_5_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110110000100"
        )
    port map (
            in0 => \N__14763\,
            in1 => \N__14840\,
            in2 => \N__14811\,
            in3 => \N__14720\,
            lcout => OPEN,
            ltout => \Lab_UT.segmentUQ_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_72_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15109\,
            in2 => \N__13798\,
            in3 => \N__19881\,
            lcout => \uu2.bitmapZ0Z_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_72C_net\,
            ce => 'H',
            sr => \N__26038\
        );

    \Lab_UT.bcd2segment3.segment_1_6_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011010"
        )
    port map (
            in0 => \N__14762\,
            in1 => \N__14839\,
            in2 => \N__14810\,
            in3 => \N__14719\,
            lcout => \Lab_UT.segment_1_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment3.segmentUQ_i_a4_1_6_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__14842\,
            in1 => \N__14796\,
            in2 => \N__14728\,
            in3 => \N__14761\,
            lcout => OPEN,
            ltout => \Lab_UT.N_65_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_168_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111010101010"
        )
    port map (
            in0 => \N__19879\,
            in1 => \N__15110\,
            in2 => \N__13795\,
            in3 => \N__13792\,
            lcout => \uu2.bitmapZ0Z_168\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_72C_net\,
            ce => 'H',
            sr => \N__26038\
        );

    \Lab_UT.bcd2segment3.segmentUQ_i_a3_4_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100001010"
        )
    port map (
            in0 => \N__14841\,
            in1 => \N__14803\,
            in2 => \N__14727\,
            in3 => \N__14764\,
            lcout => OPEN,
            ltout => \Lab_UT.N_76_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_200_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101110"
        )
    port map (
            in0 => \N__19880\,
            in1 => \N__15111\,
            in2 => \N__13786\,
            in3 => \N__13870\,
            lcout => \uu2.bitmapZ0Z_200\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_72C_net\,
            ce => 'H',
            sr => \N__26038\
        );

    \uu2.bitmap_RNIOS152_72_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011101110"
        )
    port map (
            in0 => \N__13783\,
            in1 => \N__19438\,
            in2 => \N__13777\,
            in3 => \N__14677\,
            lcout => \uu2.bitmap_RNIOS152Z0Z_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.dicLdAMtens_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__20107\,
            in1 => \N__13921\,
            in2 => \N__13939\,
            in3 => \N__17599\,
            lcout => \Lab_UT.dictrl.dicLdAMtensZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29408\,
            ce => 'H',
            sr => \N__13900\
        );

    \Lab_UT.didp.Mones_alarm.q_RNIN5N11_0_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29992\,
            in1 => \N__22765\,
            in2 => \_gnd_net_\,
            in3 => \N__19681\,
            lcout => \Lab_UT.Mone_at_0\,
            ltout => \Lab_UT.Mone_at_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment3.segmentUQ_i_a3_0_4_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13873\,
            in3 => \N__14795\,
            lcout => \Lab_UT.N_77_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Mones_alarm.q_RNITBN11_3_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28251\,
            in1 => \N__22693\,
            in2 => \_gnd_net_\,
            in3 => \N__19684\,
            lcout => \Lab_UT.Mone_at_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Mones_alarm.q_RNIP7N11_1_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__19682\,
            in1 => \N__30082\,
            in2 => \_gnd_net_\,
            in3 => \N__25780\,
            lcout => \Lab_UT.Mone_at_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Mones_alarm.q_RNIR9N11_2_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28296\,
            in1 => \N__22738\,
            in2 => \_gnd_net_\,
            in3 => \N__19683\,
            lcout => \Lab_UT.Mone_at_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Mones_subtractor.q_RNIVQVP_2_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29773\,
            in1 => \N__28297\,
            in2 => \_gnd_net_\,
            in3 => \N__26886\,
            lcout => \Lab_UT.didp.q_RNIVQVP_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__m22_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__23812\,
            in1 => \N__23976\,
            in2 => \_gnd_net_\,
            in3 => \N__15192\,
            lcout => \Lab_UT.dictrl.N_23\,
            ltout => \Lab_UT.dictrl.N_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_RNIGHD18_1_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100001010"
        )
    port map (
            in0 => \N__18007\,
            in1 => \_gnd_net_\,
            in2 => \N__13837\,
            in3 => \N__13829\,
            lcout => \Lab_UT.dictrl.nextState_RNIGHD18Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_RNIKSEU7_0_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__27783\,
            in1 => \N__21218\,
            in2 => \N__15142\,
            in3 => \N__13804\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_12_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_RNIV4IAN_1_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001010000000"
        )
    port map (
            in0 => \N__20188\,
            in1 => \N__17920\,
            in2 => \N__13951\,
            in3 => \N__17221\,
            lcout => \Lab_UT.dictrl.g0_i_a4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_RNI2P2A_2_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24964\,
            in2 => \_gnd_net_\,
            in3 => \N__23388\,
            lcout => \Lab_UT.dictrl.currState_2_RNI2P2AZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_RNI6ITB_0_2_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__23389\,
            in1 => \_gnd_net_\,
            in2 => \N__25009\,
            in3 => \N__26148\,
            lcout => \Lab_UT.dictrl.G_28_0_a5_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.dicLdAMtens_RNIDTLN4_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__13938\,
            in1 => \N__13920\,
            in2 => \_gnd_net_\,
            in3 => \N__20106\,
            lcout => \Lab_UT.ld_enable_AMtens\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__m17_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__20938\,
            in1 => \N__27782\,
            in2 => \_gnd_net_\,
            in3 => \N__27292\,
            lcout => \Lab_UT.dictrl.N_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_0_ret_10_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__14034\,
            in1 => \N__18009\,
            in2 => \N__15575\,
            in3 => \N__21044\,
            lcout => \Lab_UT.dictrl.r_dicLdMtens16_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29394\,
            ce => 'H',
            sr => \N__26063\
        );

    \Lab_UT.dictrl.currState_0_ret_17_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__21043\,
            in1 => \N__15568\,
            in2 => \N__18047\,
            in3 => \N__14035\,
            lcout => \Lab_UT.dictrl.r_dicLdMtens17_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29394\,
            ce => 'H',
            sr => \N__26063\
        );

    \Lab_UT.dictrl.r_enable1_RNO_0_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__15199\,
            in1 => \N__13909\,
            in2 => \_gnd_net_\,
            in3 => \N__17919\,
            lcout => \Lab_UT.dictrl.un1_currState_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_RNO_8_1_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__23447\,
            in1 => \N__24578\,
            in2 => \_gnd_net_\,
            in3 => \N__21536\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_10_0_N_4L6_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_RNO_3_1_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110000"
        )
    port map (
            in0 => \N__17526\,
            in1 => \N__15434\,
            in2 => \N__13903\,
            in3 => \N__21042\,
            lcout => \Lab_UT.dictrl.nextState_RNO_3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.r_enable4_RNO_0_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__17918\,
            in1 => \N__14059\,
            in2 => \N__14053\,
            in3 => \N__24863\,
            lcout => \Lab_UT.dictrl.un1_currState_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__m33_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__24862\,
            in1 => \N__17917\,
            in2 => \_gnd_net_\,
            in3 => \N__15181\,
            lcout => \Lab_UT.dictrl.N_34\,
            ltout => \Lab_UT.dictrl.N_34_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_RNIL8B7M_1_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011011111"
        )
    port map (
            in0 => \N__18008\,
            in1 => \N__24577\,
            in2 => \N__14038\,
            in3 => \N__14033\,
            lcout => \Lab_UT.dictrl.N_8ctr\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__m15_bm_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001101"
        )
    port map (
            in0 => \N__17905\,
            in1 => \N__15211\,
            in2 => \N__24861\,
            in3 => \N__14160\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.m15_bm_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_0_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14113\,
            in2 => \N__14011\,
            in3 => \N__25011\,
            lcout => \Lab_UT.dictrl.nextState_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29390\,
            ce => \N__15517\,
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_RNI1KKK6_0_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110001110100"
        )
    port map (
            in0 => \N__24815\,
            in1 => \N__18042\,
            in2 => \N__14007\,
            in3 => \N__13987\,
            lcout => \Lab_UT.dictrl.N_1609_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_3_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__13975\,
            in1 => \N__17906\,
            in2 => \N__25046\,
            in3 => \N__23785\,
            lcout => \Lab_UT.dictrl.nextState_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29390\,
            ce => \N__15517\,
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_ret_5_RNO_0_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__23784\,
            in1 => \N__18084\,
            in2 => \_gnd_net_\,
            in3 => \N__23446\,
            lcout => \Lab_UT.dictrl.currState_ret_5_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_RNI1O2A_0_1_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__23445\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17904\,
            lcout => \Lab_UT.dictrl.currState_2_RNI1O2A_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_RNI6ITB_2_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__25010\,
            in1 => \N__23444\,
            in2 => \_gnd_net_\,
            in3 => \N__26147\,
            lcout => \Lab_UT.dictrl.N_23_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__g0_16_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111110000"
        )
    port map (
            in0 => \N__27701\,
            in1 => \N__21715\,
            in2 => \N__20398\,
            in3 => \N__14194\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_14_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_RNI71NQI_1_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__18062\,
            in1 => \N__17912\,
            in2 => \N__14188\,
            in3 => \N__14185\,
            lcout => \Lab_UT.dictrl.N_1607_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__g0_8_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__20388\,
            in1 => \N__14175\,
            in2 => \_gnd_net_\,
            in3 => \N__14156\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_9_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__g0_11_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17913\,
            in2 => \N__14140\,
            in3 => \N__14131\,
            lcout => \Lab_UT.dictrl.N_10_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__g0_6_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011100001111"
        )
    port map (
            in0 => \N__27700\,
            in1 => \N__14137\,
            in2 => \N__20397\,
            in3 => \N__20295\,
            lcout => \Lab_UT.dictrl.N_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__m15_am_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101000100"
        )
    port map (
            in0 => \N__14125\,
            in1 => \N__17914\,
            in2 => \_gnd_net_\,
            in3 => \N__20283\,
            lcout => \Lab_UT.dictrl.m15_am\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_0_rep2_RNIQAFK3_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__21286\,
            in1 => \N__18375\,
            in2 => \N__20939\,
            in3 => \N__25492\,
            lcout => \Lab_UT.dictrl.N_20_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_0_rep1_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21071\,
            in2 => \_gnd_net_\,
            in3 => \N__24705\,
            lcout => \Lab_UT.dictrl.currState_0_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29384\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.decoder.de_cr_1_0_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__15669\,
            in1 => \N__15681\,
            in2 => \_gnd_net_\,
            in3 => \N__14230\,
            lcout => \Lab_UT.dictrl.de_cr_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_fast_es_RNIAJ1G_3_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__15673\,
            in1 => \N__17694\,
            in2 => \N__15685\,
            in3 => \N__15795\,
            lcout => OPEN,
            ltout => \buart.Z_rx.bitcount_fast_es_RNIAJ1GZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_RNIK0OS_0_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__15844\,
            in1 => \_gnd_net_\,
            in2 => \N__14275\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_rdy,
            ltout => \bu_rx_data_rdy_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_fast_RNIC98T_0_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14272\,
            in3 => \N__14509\,
            lcout => \Lab_UT.dictrl.N_5_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__g1_0_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__24357\,
            in1 => \N__28979\,
            in2 => \_gnd_net_\,
            in3 => \N__24414\,
            lcout => \Lab_UT.dictrl.g1_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.decoder.g0_3_1_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__28978\,
            in1 => \N__28606\,
            in2 => \_gnd_net_\,
            in3 => \N__24358\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__g0_1_1_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110011001100"
        )
    port map (
            in0 => \N__24207\,
            in1 => \N__21246\,
            in2 => \N__14242\,
            in3 => \N__27712\,
            lcout => \Lab_UT.dictrl.g0_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_fast_0_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__28812\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_fast_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29381\,
            ce => \N__25429\,
            sr => \N__26091\
        );

    \Lab_UT.dictrl.decoder.de_num_1_2_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__14328\,
            in1 => \N__14304\,
            in2 => \N__14362\,
            in3 => \N__14313\,
            lcout => \Lab_UT.dictrl.de_num_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.decoder.g0_0_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__21895\,
            in1 => \N__17617\,
            in2 => \N__15496\,
            in3 => \N__14361\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.decoder.g0_5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.decoder.g0_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14338\,
            in1 => \N__14320\,
            in2 => \N__14350\,
            in3 => \N__17649\,
            lcout => \Lab_UT.dictrl.de_cr_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.decoder.g0_3_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__14314\,
            in1 => \N__20839\,
            in2 => \N__15843\,
            in3 => \N__15796\,
            lcout => \Lab_UT.dictrl.decoder.g0_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.decoder.g0_4_LC_5_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__14329\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14305\,
            lcout => \Lab_UT.dictrl.decoder.g0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_fast_4_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24417\,
            lcout => bu_rx_data_fast_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29376\,
            ce => \N__25426\,
            sr => \N__26094\
        );

    \buart.Z_rx.shifter_fast_5_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__24271\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_fast_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29376\,
            ce => \N__25426\,
            sr => \N__26094\
        );

    \buart.Z_rx.shifter_5_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24270\,
            lcout => bu_rx_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29376\,
            ce => \N__25426\,
            sr => \N__26094\
        );

    \buart.Z_rx.hh_RNIJ3K62_0_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__15636\,
            in1 => \_gnd_net_\,
            in2 => \N__14296\,
            in3 => \N__21872\,
            lcout => \buart.Z_rx.startbit\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.decoder.g0_9_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__21764\,
            in1 => \N__21935\,
            in2 => \N__21995\,
            in3 => \N__17698\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.decoder.g0Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.decoder.g0_2_LC_5_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15658\,
            in1 => \N__14443\,
            in2 => \N__14512\,
            in3 => \N__18171\,
            lcout => \Lab_UT.dictrl.de_littleA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__g1_4_1_LC_5_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111111111111"
        )
    port map (
            in0 => \N__21986\,
            in1 => \_gnd_net_\,
            in2 => \N__14508\,
            in3 => \N__21696\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g1_4_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__g1_4_LC_5_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__24440\,
            in1 => \N__21765\,
            in2 => \N__14467\,
            in3 => \N__24356\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__g0_10_LC_5_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100010111011"
        )
    port map (
            in0 => \N__24003\,
            in1 => \N__14464\,
            in2 => \N__14458\,
            in3 => \N__27725\,
            lcout => \Lab_UT.dictrl.N_17_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.decoder.g0_7_LC_5_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__21394\,
            in1 => \N__25260\,
            in2 => \_gnd_net_\,
            in3 => \N__21697\,
            lcout => \Lab_UT.dictrl.decoder.g0_5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__m7_sx_LC_5_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__21763\,
            in1 => \N__21695\,
            in2 => \N__24012\,
            in3 => \N__21393\,
            lcout => \Lab_UT.dictrl.m7_sx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_0_LC_5_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15922\,
            in2 => \_gnd_net_\,
            in3 => \N__14414\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29371\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_RNI3O55_3_LC_5_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__14427\,
            in1 => \N__14413\,
            in2 => \_gnd_net_\,
            in3 => \N__14395\,
            lcout => \buart.Z_rx.ser_clk\,
            ltout => \buart.Z_rx.ser_clk_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_4_LC_5_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000100"
        )
    port map (
            in0 => \N__15921\,
            in1 => \N__14389\,
            in2 => \N__14383\,
            in3 => \N__14379\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29371\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_RNIGD8S2_1_LC_5_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__15637\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27729\,
            lcout => \buart.Z_rx.N_27_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_0_LC_6_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010011001"
        )
    port map (
            in0 => \N__19172\,
            in1 => \N__19218\,
            in2 => \_gnd_net_\,
            in3 => \N__20433\,
            lcout => \resetGen.reset_countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29437\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_RNO_0_4_LC_6_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18937\,
            in2 => \_gnd_net_\,
            in3 => \N__19144\,
            lcout => OPEN,
            ltout => \resetGen.reset_count_2_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_4_LC_6_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011101100"
        )
    port map (
            in0 => \N__19204\,
            in1 => \N__19171\,
            in2 => \N__14566\,
            in3 => \N__20434\,
            lcout => \resetGen.reset_countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29437\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_1_LC_6_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__19035\,
            in1 => \N__18771\,
            in2 => \_gnd_net_\,
            in3 => \N__14917\,
            lcout => \uu2.mem0.w_addr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_3_LC_6_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__18772\,
            in1 => \N__22460\,
            in2 => \_gnd_net_\,
            in3 => \N__16505\,
            lcout => \uu2.mem0.w_addr_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_w_addr_user.counter_gen_label_6__un426_ci_3_LC_6_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__22461\,
            in1 => \_gnd_net_\,
            in2 => \N__22492\,
            in3 => \_gnd_net_\,
            lcout => \uu2.un426_ci_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_4_LC_6_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__18773\,
            in1 => \N__22488\,
            in2 => \_gnd_net_\,
            in3 => \N__16543\,
            lcout => \uu2.mem0.w_addr_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_5_LC_6_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22351\,
            in1 => \N__16446\,
            in2 => \_gnd_net_\,
            in3 => \N__18774\,
            lcout => \uu2.mem0.w_addr_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIGEPH1_4_LC_6_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110010000000"
        )
    port map (
            in0 => \N__16256\,
            in1 => \N__16504\,
            in2 => \N__16121\,
            in3 => \N__14909\,
            lcout => \uu2.bitmap_pmux_sn_N_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNI6RO21_162_LC_6_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__14620\,
            in1 => \N__16253\,
            in2 => \_gnd_net_\,
            in3 => \N__14938\,
            lcout => OPEN,
            ltout => \uu2.N_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNIELSJ2_111_LC_6_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14596\,
            in2 => \N__14611\,
            in3 => \N__14602\,
            lcout => \uu2.bitmap_RNIELSJ2Z0Z_111\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIM0T61_2_LC_6_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000010001"
        )
    port map (
            in0 => \N__14907\,
            in1 => \N__16254\,
            in2 => \_gnd_net_\,
            in3 => \N__16103\,
            lcout => \uu2.bitmap_pmux_sn_N_54_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_111_LC_6_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26800\,
            lcout => \uu2.bitmapZ0Z_111\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_111C_net\,
            ce => 'H',
            sr => \N__26046\
        );

    \uu2.w_addr_displaying_RNI8NSO_4_LC_6_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16498\,
            in2 => \_gnd_net_\,
            in3 => \N__16104\,
            lcout => \uu2.bitmap_pmux_sn_N_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI8NSO_2_LC_6_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__16255\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14908\,
            lcout => \uu2.N_39\,
            ltout => \uu2.N_39_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_w_addr_displaying.result_1_0_o2_4_LC_6_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19496\,
            in2 => \N__14569\,
            in3 => \N__16108\,
            lcout => \uu2.N_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_nesr_3_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__16120\,
            in1 => \N__14906\,
            in2 => \N__19497\,
            in3 => \N__16271\,
            lcout => \uu2.w_addr_displayingZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_nesr_3C_net\,
            ce => \N__16303\,
            sr => \N__26044\
        );

    \uu2.w_addr_displaying_nesr_1_LC_6_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19483\,
            in2 => \_gnd_net_\,
            in3 => \N__16119\,
            lcout => \uu2.w_addr_displayingZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_nesr_3C_net\,
            ce => \N__16303\,
            sr => \N__26044\
        );

    \uu2.w_addr_displaying_nesr_7_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100110101010"
        )
    port map (
            in0 => \N__16778\,
            in1 => \N__16461\,
            in2 => \N__16374\,
            in3 => \N__16441\,
            lcout => \uu2.w_addr_displayingZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_nesr_3C_net\,
            ce => \N__16303\,
            sr => \N__26044\
        );

    \uu2.w_addr_displaying_ness_6_LC_6_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101011010101"
        )
    port map (
            in0 => \N__16440\,
            in1 => \N__16777\,
            in2 => \N__16639\,
            in3 => \N__14671\,
            lcout => \uu2.w_addr_displayingZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_nesr_3C_net\,
            ce => \N__16303\,
            sr => \N__26044\
        );

    \CONSTANT_ONE_LUT4_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNI35M31_84_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010100101111"
        )
    port map (
            in0 => \N__16757\,
            in1 => \N__14653\,
            in2 => \N__19459\,
            in3 => \N__16900\,
            lcout => \uu2.bitmap_pmux_24_am_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_87_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__19882\,
            in1 => \N__16294\,
            in2 => \_gnd_net_\,
            in3 => \N__20170\,
            lcout => \uu2.bitmapZ0Z_87\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_87C_net\,
            ce => 'H',
            sr => \N__26042\
        );

    \uu2.bitmap_314_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__19543\,
            in1 => \N__19883\,
            in2 => \_gnd_net_\,
            in3 => \N__19096\,
            lcout => \uu2.bitmapZ0Z_314\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_87C_net\,
            ce => 'H',
            sr => \N__26042\
        );

    \uu2.bitmap_RNIVKR41_180_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16678\,
            in2 => \N__16272\,
            in3 => \N__14640\,
            lcout => OPEN,
            ltout => \uu2.N_386_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_nesr_RNI1JET2_7_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__16756\,
            in1 => \N__16250\,
            in2 => \N__14647\,
            in3 => \N__16558\,
            lcout => OPEN,
            ltout => \uu2.w_addr_displaying_nesr_RNI1JET2Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNIMAS54_314_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100101111"
        )
    port map (
            in0 => \N__16252\,
            in1 => \N__16110\,
            in2 => \N__14644\,
            in3 => \N__14641\,
            lcout => \uu2.bitmap_pmux_23_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIAGTK1_2_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100000110"
        )
    port map (
            in0 => \N__14898\,
            in1 => \N__16109\,
            in2 => \N__16779\,
            in3 => \N__16251\,
            lcout => \uu2.bitmap_pmux_sn_N_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_2_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__19473\,
            in1 => \N__14899\,
            in2 => \N__16336\,
            in3 => \N__16111\,
            lcout => \uu2.w_addr_displayingZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_87C_net\,
            ce => 'H',
            sr => \N__26042\
        );

    \Lab_UT.didp.Mones_alarm.q_RNI83T64_1_1_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010010010"
        )
    port map (
            in0 => \N__14835\,
            in1 => \N__14804\,
            in2 => \N__14765\,
            in3 => \N__14715\,
            lcout => \Lab_UT.L3_segment3_0_i_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Mones_alarm.q_RNI83T64_1_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011011011"
        )
    port map (
            in0 => \N__14716\,
            in1 => \N__14754\,
            in2 => \N__14812\,
            in3 => \N__14836\,
            lcout => \Lab_UT.L3_segment3_0_i_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Mones_alarm.q_RNI83T64_0_1_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111010111111"
        )
    port map (
            in0 => \N__14837\,
            in1 => \N__14808\,
            in2 => \N__14766\,
            in3 => \N__14717\,
            lcout => OPEN,
            ltout => \Lab_UT.L3_segment3_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_203_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15107\,
            in2 => \N__14845\,
            in3 => \N__19893\,
            lcout => \uu2.bitmapZ0Z_203\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_203C_net\,
            ce => 'H',
            sr => \N__26040\
        );

    \Lab_UT.didp.Mones_alarm.q_RNI83T64_2_1_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011110011111"
        )
    port map (
            in0 => \N__14838\,
            in1 => \N__14809\,
            in2 => \N__14767\,
            in3 => \N__14718\,
            lcout => OPEN,
            ltout => \Lab_UT.L3_segment3_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_75_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15108\,
            in2 => \N__14692\,
            in3 => \N__19894\,
            lcout => \uu2.bitmapZ0Z_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_203C_net\,
            ce => 'H',
            sr => \N__26040\
        );

    \uu2.bitmap_RNI99H91_75_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000001011111"
        )
    port map (
            in0 => \N__14689\,
            in1 => \N__14683\,
            in2 => \N__19458\,
            in3 => \N__16780\,
            lcout => \uu2.bitmap_pmux_24_bm_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_0_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__16332\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19425\,
            lcout => \uu2.w_addr_displayingZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_203C_net\,
            ce => 'H',
            sr => \N__26040\
        );

    \Lab_UT.bcd2segment4.segmentUQ_i_a3_4_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000101110"
        )
    port map (
            in0 => \N__17041\,
            in1 => \N__19604\,
            in2 => \N__17001\,
            in3 => \N__16940\,
            lcout => OPEN,
            ltout => \Lab_UT.N_76_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_194_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000100"
        )
    port map (
            in0 => \N__16948\,
            in1 => \N__15055\,
            in2 => \N__14983\,
            in3 => \N__19896\,
            lcout => \uu2.bitmapZ0Z_194\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_194C_net\,
            ce => 'H',
            sr => \N__26037\
        );

    \Lab_UT.didp.Mtens_alarm.q_RNIGGJ64_2_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000010000110"
        )
    port map (
            in0 => \N__17040\,
            in1 => \N__19603\,
            in2 => \N__17000\,
            in3 => \N__16939\,
            lcout => \Lab_UT.L3_segment4_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Mtens_alarm.q_RNIGGJ64_0_2_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011100011111"
        )
    port map (
            in0 => \N__16941\,
            in1 => \N__16994\,
            in2 => \N__19609\,
            in3 => \N__17042\,
            lcout => OPEN,
            ltout => \Lab_UT.L3_segment4_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_69_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15039\,
            in2 => \N__14968\,
            in3 => \N__19820\,
            lcout => \uu2.bitmapZ0Z_69\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_194C_net\,
            ce => 'H',
            sr => \N__26037\
        );

    \uu2.bitmap_34_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001010"
        )
    port map (
            in0 => \N__15038\,
            in1 => \_gnd_net_\,
            in2 => \N__19875\,
            in3 => \N__14956\,
            lcout => \uu2.bitmapZ0Z_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_194C_net\,
            ce => 'H',
            sr => \N__26037\
        );

    \Lab_UT.bcd2segment4.segment_1_6_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111100"
        )
    port map (
            in0 => \N__17043\,
            in1 => \N__19608\,
            in2 => \N__17002\,
            in3 => \N__16942\,
            lcout => OPEN,
            ltout => \Lab_UT.segment_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_162_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011101100"
        )
    port map (
            in0 => \N__15040\,
            in1 => \N__19895\,
            in2 => \N__14941\,
            in3 => \N__16882\,
            lcout => \uu2.bitmapZ0Z_162\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_194C_net\,
            ce => 'H',
            sr => \N__26037\
        );

    \Lab_UT.dictrl.nextState_RNI6VQ05_2_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010100000"
        )
    port map (
            in0 => \N__18130\,
            in1 => \N__15537\,
            in2 => \N__20857\,
            in3 => \N__23436\,
            lcout => \Lab_UT.dictrl.N_1614_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_0_ret_21_RNIUL8L_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__18013\,
            in1 => \N__23813\,
            in2 => \_gnd_net_\,
            in3 => \N__24006\,
            lcout => \Lab_UT.dictrl.N_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.r_enable1_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111001010"
        )
    port map (
            in0 => \N__15133\,
            in1 => \N__15127\,
            in2 => \N__23457\,
            in3 => \N__20200\,
            lcout => \Lab_UT.dictrl.r_enableZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29393\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.r_enable1_RNI7DR61_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__15126\,
            in1 => \N__24168\,
            in2 => \N__23176\,
            in3 => \N__23654\,
            lcout => \Lab_UT.dictrl.enableSeg1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.r_enable3_RNI9DR61_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__23655\,
            in1 => \N__15072\,
            in2 => \N__24176\,
            in3 => \N__23174\,
            lcout => \Lab_UT.dictrl.enableSeg3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.r_enable3_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__23437\,
            in1 => \N__19695\,
            in2 => \N__15076\,
            in3 => \N__21307\,
            lcout => \Lab_UT.dictrl.r_enableZ0Z3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29393\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.r_enable4_RNIADR61_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__23656\,
            in1 => \N__15000\,
            in2 => \N__24177\,
            in3 => \N__23175\,
            lcout => \Lab_UT.dictrl.enableSeg4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.r_enable4_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010110001"
        )
    port map (
            in0 => \N__23438\,
            in1 => \N__19696\,
            in2 => \N__15004\,
            in3 => \N__15013\,
            lcout => \Lab_UT.dictrl.r_enableZ0Z4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29393\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_RNI19TAN_1_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__14992\,
            in1 => \N__17911\,
            in2 => \_gnd_net_\,
            in3 => \N__17230\,
            lcout => \Lab_UT.dictrl.g1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_RNI421C4_0_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__27285\,
            in1 => \N__21250\,
            in2 => \N__27810\,
            in3 => \N__17442\,
            lcout => \Lab_UT.dictrl.N_17_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__g0_19_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__17629\,
            in1 => \N__27777\,
            in2 => \N__21264\,
            in3 => \N__27284\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_36_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_RNIBR9BG_1_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17443\,
            in2 => \N__15205\,
            in3 => \N__17452\,
            lcout => \Lab_UT.dictrl.nextStateZ0Z_3\,
            ltout => \Lab_UT.dictrl.nextStateZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_0_ret_26_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24682\,
            in2 => \N__15202\,
            in3 => \N__21072\,
            lcout => \Lab_UT.dictrl.r_dicLdMtens21_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29388\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_0_ret_25_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__17546\,
            in1 => \N__15474\,
            in2 => \N__17356\,
            in3 => \N__15385\,
            lcout => \Lab_UT.dictrl.r_dicLdMtens22_i_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29388\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_0_ret_27_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__15475\,
            in1 => \N__17355\,
            in2 => \N__17335\,
            in3 => \N__17547\,
            lcout => \Lab_UT.dictrl.r_dicLdMtens20_i_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29388\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__m32_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000001110101"
        )
    port map (
            in0 => \N__23816\,
            in1 => \N__24481\,
            in2 => \N__21265\,
            in3 => \N__15193\,
            lcout => \Lab_UT.dictrl.N_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_RNIDED951_2_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011001101"
        )
    port map (
            in0 => \N__23453\,
            in1 => \N__15175\,
            in2 => \N__25047\,
            in3 => \N__15169\,
            lcout => \Lab_UT.dictrl.nextStateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_RNID73K33_1_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011101111111"
        )
    port map (
            in0 => \N__21035\,
            in1 => \N__15163\,
            in2 => \N__21609\,
            in3 => \N__20751\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_0_ret_29_RNIOSJNC6_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__23454\,
            in1 => \N__24677\,
            in2 => \N__15286\,
            in3 => \N__17128\,
            lcout => \Lab_UT.dictrl.g0_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_RNO_9_1_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__24678\,
            in1 => \N__23455\,
            in2 => \_gnd_net_\,
            in3 => \N__20668\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.nextState_RNO_9Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_RNO_4_1_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__15279\,
            in1 => \N__15244\,
            in2 => \N__15283\,
            in3 => \N__17122\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.nextState_RNO_4Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_RNO_1_1_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110000"
        )
    port map (
            in0 => \N__15280\,
            in1 => \N__15238\,
            in2 => \N__15262\,
            in3 => \N__15259\,
            lcout => \Lab_UT.dictrl.g0_i_o4_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_RNO_11_1_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21568\,
            in2 => \N__20795\,
            in3 => \N__21036\,
            lcout => \Lab_UT.dictrl.N_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_RNO_5_1_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000110000"
        )
    port map (
            in0 => \N__17532\,
            in1 => \N__20755\,
            in2 => \N__21610\,
            in3 => \N__15484\,
            lcout => \Lab_UT.dictrl.N_18_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__g0_23_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001011111010"
        )
    port map (
            in0 => \N__21259\,
            in1 => \N__27710\,
            in2 => \N__18343\,
            in3 => \N__27299\,
            lcout => \Lab_UT.dictrl.N_13_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__g1_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__23831\,
            in1 => \N__24309\,
            in2 => \N__15232\,
            in3 => \N__28602\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g1_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__g0_22_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011101110"
        )
    port map (
            in0 => \N__15223\,
            in1 => \N__23832\,
            in2 => \N__15214\,
            in3 => \N__27711\,
            lcout => \Lab_UT.dictrl.N_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_0_ret_28_RNO_0_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__17351\,
            in1 => \N__17553\,
            in2 => \N__17331\,
            in3 => \N__15481\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.r_dicLdMtens20_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_0_ret_28_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000001100"
        )
    port map (
            in0 => \N__15409\,
            in1 => \N__17488\,
            in2 => \N__15487\,
            in3 => \N__15358\,
            lcout => \Lab_UT.dictrl.r_Sone_init17_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29379\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_RNIFGT042_0_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17552\,
            in2 => \_gnd_net_\,
            in3 => \N__15480\,
            lcout => \Lab_UT.dictrl.r_dicLdMtens22_2_reti\,
            ltout => \Lab_UT.dictrl.r_dicLdMtens22_2_reti_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_0_ret_29_RNIDFRSEE_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100000000"
        )
    port map (
            in0 => \N__15403\,
            in1 => \N__15357\,
            in2 => \N__15394\,
            in3 => \N__15391\,
            lcout => \Lab_UT.dictrl.currState_0_ret_29_RNIDFRSEEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_0_ret_21_RNIPJM6D1_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__17350\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15384\,
            lcout => \Lab_UT.dictrl.r_dicLdMtens22_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__m27_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__15297\,
            in1 => \N__21267\,
            in2 => \_gnd_net_\,
            in3 => \N__24874\,
            lcout => \Lab_UT.dictrl.N_41_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_RNIN9NP3_7_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111111111111"
        )
    port map (
            in0 => \N__25397\,
            in1 => \N__21290\,
            in2 => \N__18376\,
            in3 => \N__25478\,
            lcout => \N_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__m29_LC_6_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011110101111"
        )
    port map (
            in0 => \N__23798\,
            in1 => \N__17099\,
            in2 => \N__15337\,
            in3 => \N__21266\,
            lcout => \Lab_UT.dictrl.N_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.decoder.de_littleA_LC_6_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__25398\,
            in1 => \N__17473\,
            in2 => \N__24208\,
            in3 => \N__21291\,
            lcout => \Lab_UT.dictrl.de_littleA\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.decoder.de_cr_1_LC_6_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__18224\,
            in1 => \N__18179\,
            in2 => \_gnd_net_\,
            in3 => \N__17650\,
            lcout => \Lab_UT_dictrl_decoder_de_cr_1\,
            ltout => \Lab_UT_dictrl_decoder_de_cr_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.decoder.de_cr_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__18371\,
            in1 => \N__25394\,
            in2 => \N__15598\,
            in3 => \N__25477\,
            lcout => \Lab_UT.dictrl.de_cr\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__m30_LC_6_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__17928\,
            in1 => \N__15595\,
            in2 => \_gnd_net_\,
            in3 => \N__15589\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_2_LC_6_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15582\,
            in2 => \N__15544\,
            in3 => \N__25040\,
            lcout => \Lab_UT.dictrl.nextState_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29374\,
            ce => \N__15513\,
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_fast_es_2_LC_6_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0010011101110010"
        )
    port map (
            in0 => \N__15977\,
            in1 => \N__15931\,
            in2 => \N__15745\,
            in3 => \N__18236\,
            lcout => \buart__rx_bitcount_fast_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29372\,
            ce => \N__15870\,
            sr => \N__26095\
        );

    \buart.Z_rx.bitcount_es_2_LC_6_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0001110100101110"
        )
    port map (
            in0 => \N__18235\,
            in1 => \N__15974\,
            in2 => \N__15941\,
            in3 => \N__15740\,
            lcout => \buart__rx_bitcount_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29372\,
            ce => \N__15870\,
            sr => \N__26095\
        );

    \buart.Z_rx.bitcount_2_rep1_es_LC_6_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0010011101110010"
        )
    port map (
            in0 => \N__15972\,
            in1 => \N__15928\,
            in2 => \N__15744\,
            in3 => \N__18234\,
            lcout => \buart__rx_bitcount_2_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29372\,
            ce => \N__15870\,
            sr => \N__26095\
        );

    \buart.Z_rx.bitcount_es_1_LC_6_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0100011101110100"
        )
    port map (
            in0 => \N__15927\,
            in1 => \N__15973\,
            in2 => \N__15760\,
            in3 => \N__15803\,
            lcout => \buart__rx_bitcount_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29372\,
            ce => \N__15870\,
            sr => \N__26095\
        );

    \buart.Z_rx.bitcount_es_4_LC_6_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0010011101110010"
        )
    port map (
            in0 => \N__15976\,
            in1 => \N__15930\,
            in2 => \N__15700\,
            in3 => \N__18319\,
            lcout => \buart__rx_bitcount_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29372\,
            ce => \N__15870\,
            sr => \N__26095\
        );

    \buart.Z_rx.bitcount_fast_es_4_LC_6_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0001110100101110"
        )
    port map (
            in0 => \N__18318\,
            in1 => \N__15979\,
            in2 => \N__15943\,
            in3 => \N__15699\,
            lcout => \buart__rx_bitcount_fast_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29372\,
            ce => \N__15870\,
            sr => \N__26095\
        );

    \buart.Z_rx.bitcount_es_3_LC_6_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0010011101110010"
        )
    port map (
            in0 => \N__15975\,
            in1 => \N__15929\,
            in2 => \N__15721\,
            in3 => \N__18278\,
            lcout => \buart__rx_bitcount_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29372\,
            ce => \N__15870\,
            sr => \N__26095\
        );

    \buart.Z_rx.bitcount_fast_es_3_LC_6_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0001110100101110"
        )
    port map (
            in0 => \N__18279\,
            in1 => \N__15978\,
            in2 => \N__15942\,
            in3 => \N__15720\,
            lcout => \buart__rx_bitcount_fast_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29372\,
            ce => \N__15870\,
            sr => \N__26095\
        );

    \Lab_UT.dictrl.decoder.g0_8_LC_6_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__18269\,
            in1 => \N__21837\,
            in2 => \N__18321\,
            in3 => \N__21351\,
            lcout => \Lab_UT.dictrl.decoder.g0_6_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_RNIIVPI1_1_LC_6_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__18232\,
            in1 => \N__18270\,
            in2 => \N__15804\,
            in3 => \N__18317\,
            lcout => OPEN,
            ltout => \buart.Z_rx.un1_sample_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_RNIV4M42_0_LC_6_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__15837\,
            in1 => \_gnd_net_\,
            in2 => \N__15652\,
            in3 => \N__15619\,
            lcout => \buart.Z_rx.sample\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_RNILRCP_0_LC_6_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15835\,
            in2 => \_gnd_net_\,
            in3 => \N__15793\,
            lcout => \buart__rx_valid_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_RNIOUCP_0_LC_6_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__15836\,
            in1 => \_gnd_net_\,
            in2 => \N__18322\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \buart.Z_rx.idle_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_RNISCGV1_1_LC_6_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18233\,
            in1 => \N__18271\,
            in2 => \N__15640\,
            in3 => \N__15794\,
            lcout => \buart.Z_rx.idle\,
            ltout => \buart.Z_rx.idle_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_fast_sbtinv_3_LC_6_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101110"
        )
    port map (
            in0 => \N__15919\,
            in1 => \N__15620\,
            in2 => \N__15601\,
            in3 => \N__27781\,
            lcout => \buart.Z_rx.bitcounte_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_0_LC_6_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0010011101110010"
        )
    port map (
            in0 => \N__15954\,
            in1 => \N__15920\,
            in2 => \N__28356\,
            in3 => \N__15838\,
            lcout => \buart__rx_bitcount_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29370\,
            ce => \N__15871\,
            sr => \N__26096\
        );

    \buart.Z_rx.bitcount_cry_c_0_LC_6_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15842\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_16_0_\,
            carryout => \buart.Z_rx.bitcount_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_6_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15805\,
            in2 => \_gnd_net_\,
            in3 => \N__15748\,
            lcout => \buart.Z_rx.bitcount_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.bitcount_cry_0\,
            carryout => \buart.Z_rx.bitcount_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_6_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18238\,
            in2 => \_gnd_net_\,
            in3 => \N__15724\,
            lcout => \buart.Z_rx.bitcount_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.bitcount_cry_1\,
            carryout => \buart.Z_rx.bitcount_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_6_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18280\,
            in2 => \_gnd_net_\,
            in3 => \N__15706\,
            lcout => \buart.Z_rx.bitcount_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.bitcount_cry_2\,
            carryout => \buart.Z_rx.bitcount_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_3_THRU_LUT4_0_LC_6_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15703\,
            lcout => \buart.Z_rx.bitcount_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.decoder.g0_3_0_LC_6_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__28974\,
            in1 => \N__18237\,
            in2 => \_gnd_net_\,
            in3 => \N__28601\,
            lcout => \Lab_UT.dictrl.decoder.g0_3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.uu0.l_count_18_LC_7_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__18460\,
            in1 => \N__22071\,
            in2 => \_gnd_net_\,
            in3 => \N__23248\,
            lcout => \Lab_UT.uu0.l_countZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29463\,
            ce => \N__22174\,
            sr => \N__26099\
        );

    \Lab_UT.uu0.l_count_13_LC_7_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__18602\,
            in1 => \N__16029\,
            in2 => \N__15988\,
            in3 => \N__23247\,
            lcout => \Lab_UT.uu0.l_countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29463\,
            ce => \N__22174\,
            sr => \N__26099\
        );

    \Lab_UT.uu0.l_count_2_LC_7_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21793\,
            in2 => \_gnd_net_\,
            in3 => \N__22241\,
            lcout => \Lab_UT.uu0.l_countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29463\,
            ce => \N__22174\,
            sr => \N__26099\
        );

    \Lab_UT.uu0.l_count_RNIFRMN_3_LC_7_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__18450\,
            in1 => \N__18500\,
            in2 => \N__18487\,
            in3 => \N__22264\,
            lcout => \Lab_UT.uu0.un4_l_count_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.uu0.l_count_12_LC_7_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001001000100010"
        )
    port map (
            in0 => \N__16005\,
            in1 => \N__23240\,
            in2 => \N__18694\,
            in3 => \N__18604\,
            lcout => \Lab_UT.uu0.l_countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29456\,
            ce => \N__22172\,
            sr => \N__26098\
        );

    \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_7_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__18558\,
            in1 => \N__18452\,
            in2 => \_gnd_net_\,
            in3 => \N__18430\,
            lcout => OPEN,
            ltout => \Lab_UT.uu0.un143_ci_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.uu0.l_count_11_LC_7_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001001000100010"
        )
    port map (
            in0 => \N__22560\,
            in1 => \N__23239\,
            in2 => \N__16015\,
            in3 => \N__18603\,
            lcout => \Lab_UT.uu0.l_countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29456\,
            ce => \N__22172\,
            sr => \N__26098\
        );

    \Lab_UT.uu0.l_count_9_LC_7_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__18559\,
            in1 => \_gnd_net_\,
            in2 => \N__18610\,
            in3 => \N__18453\,
            lcout => \Lab_UT.uu0.l_countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29456\,
            ce => \N__22172\,
            sr => \N__26098\
        );

    \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_7_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18451\,
            in1 => \N__18429\,
            in2 => \N__22561\,
            in3 => \N__18557\,
            lcout => \Lab_UT.uu0.un154_ci_9\,
            ltout => \Lab_UT.uu0.un154_ci_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_7_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16012\,
            in3 => \N__16004\,
            lcout => \Lab_UT.uu0.un165_ci_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_RNI1VU6_3_LC_7_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__22487\,
            in1 => \N__18991\,
            in2 => \N__16155\,
            in3 => \N__19049\,
            lcout => \uu2.un3_w_addr_user_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_RNI7UV5_8_LC_7_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__22459\,
            in1 => \N__16172\,
            in2 => \_gnd_net_\,
            in3 => \N__18962\,
            lcout => OPEN,
            ltout => \uu2.un3_w_addr_user_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_RNIINVH_2_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__22352\,
            in1 => \N__19030\,
            in2 => \N__16285\,
            in3 => \N__16282\,
            lcout => \uu2.un3_w_addr_user\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_3_LC_7_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__19050\,
            in1 => \N__18993\,
            in2 => \N__19036\,
            in3 => \N__18963\,
            lcout => \uu2.w_addr_userZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_nesr_3C_net\,
            ce => \N__18535\,
            sr => \N__22322\
        );

    \uu2.mem0.ram512X8_inst_RNO_2_LC_7_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__18992\,
            in1 => \N__18749\,
            in2 => \_gnd_net_\,
            in3 => \N__16276\,
            lcout => \uu2.mem0.w_addr_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_w_addr_user.counter_gen_label_8__un448_ci_0_LC_7_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22353\,
            in2 => \_gnd_net_\,
            in3 => \N__16150\,
            lcout => OPEN,
            ltout => \uu2.vbuf_w_addr_user.un448_ci_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_8_LC_7_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__16173\,
            in1 => \N__22370\,
            in2 => \N__16180\,
            in3 => \N__22399\,
            lcout => \uu2.w_addr_userZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_nesr_3C_net\,
            ce => \N__18535\,
            sr => \N__22322\
        );

    \uu2.w_addr_user_nesr_7_LC_7_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__22398\,
            in1 => \N__22354\,
            in2 => \N__22374\,
            in3 => \N__16151\,
            lcout => \uu2.w_addr_userZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_nesr_3C_net\,
            ce => \N__18535\,
            sr => \N__22322\
        );

    \uu2.w_addr_displaying_RNIHGM43_8_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__16118\,
            in1 => \N__16388\,
            in2 => \N__16052\,
            in3 => \N__16616\,
            lcout => \uu2.N_71\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_8_LC_7_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011000110"
        )
    port map (
            in0 => \N__16331\,
            in1 => \N__16618\,
            in2 => \N__16397\,
            in3 => \N__16364\,
            lcout => \uu2.w_addr_displayingZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_8C_net\,
            ce => 'H',
            sr => \N__26049\
        );

    \uu2.w_addr_displaying_4_LC_7_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101101000100"
        )
    port map (
            in0 => \N__16362\,
            in1 => \N__16329\,
            in2 => \_gnd_net_\,
            in3 => \N__16500\,
            lcout => \uu2.w_addr_displayingZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_8C_net\,
            ce => 'H',
            sr => \N__26049\
        );

    \uu2.w_addr_displaying_5_LC_7_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001111000"
        )
    port map (
            in0 => \N__16330\,
            in1 => \N__16506\,
            in2 => \N__16544\,
            in3 => \N__16363\,
            lcout => \uu2.w_addr_displayingZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_8C_net\,
            ce => 'H',
            sr => \N__26049\
        );

    \uu2.w_addr_displaying_RNILSOL_5_LC_7_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16533\,
            in2 => \_gnd_net_\,
            in3 => \N__16499\,
            lcout => \uu2.N_41\,
            ltout => \uu2.N_41_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_ness_RNITTSI1_6_LC_7_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16433\,
            in2 => \N__16402\,
            in3 => \N__16771\,
            lcout => \uu2.N_43\,
            ltout => \uu2.N_43_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIFCPV4_8_LC_7_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011100110011"
        )
    port map (
            in0 => \N__16361\,
            in1 => \N__18748\,
            in2 => \N__16339\,
            in3 => \N__16617\,
            lcout => \uu2.w_addr_displaying_RNIFCPV4Z0Z_8\,
            ltout => \uu2.w_addr_displaying_RNIFCPV4Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIJ5K15_8_LC_7_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16306\,
            in3 => \N__26146\,
            lcout => \uu2.N_36_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Stens_alarm.q_RNI0QLC5_2_1_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101110110111"
        )
    port map (
            in0 => \N__20044\,
            in1 => \N__19938\,
            in2 => \N__20008\,
            in3 => \N__20074\,
            lcout => \Lab_UT.L3_segment2_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Stens_alarm.q_RNI0QLC5_1_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101011100111"
        )
    port map (
            in0 => \N__20077\,
            in1 => \N__20007\,
            in2 => \N__19951\,
            in3 => \N__20047\,
            lcout => OPEN,
            ltout => \Lab_UT.L3_segment2_0_i_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_308_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101010101010"
        )
    port map (
            in0 => \N__19849\,
            in1 => \_gnd_net_\,
            in2 => \N__16288\,
            in3 => \N__20168\,
            lcout => \uu2.bitmapZ0Z_308\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_308C_net\,
            ce => 'H',
            sr => \N__26047\
        );

    \Lab_UT.didp.Stens_alarm.q_RNI0QLC5_0_1_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111100111101"
        )
    port map (
            in0 => \N__20075\,
            in1 => \N__20005\,
            in2 => \N__19949\,
            in3 => \N__20045\,
            lcout => OPEN,
            ltout => \Lab_UT.L3_segment2_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_215_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__19848\,
            in1 => \_gnd_net_\,
            in2 => \N__16672\,
            in3 => \N__20167\,
            lcout => \uu2.bitmapZ0Z_215\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_308C_net\,
            ce => 'H',
            sr => \N__26047\
        );

    \Lab_UT.didp.Stens_alarm.q_RNI0QLC5_1_1_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100100010000"
        )
    port map (
            in0 => \N__20076\,
            in1 => \N__20006\,
            in2 => \N__19950\,
            in3 => \N__20046\,
            lcout => OPEN,
            ltout => \Lab_UT.L3_segment2_0_i_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_52_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110101010"
        )
    port map (
            in0 => \N__19850\,
            in1 => \_gnd_net_\,
            in2 => \N__16654\,
            in3 => \N__20169\,
            lcout => \uu2.bitmapZ0Z_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_308C_net\,
            ce => 'H',
            sr => \N__26047\
        );

    \uu2.bitmap_RNIU2IS_52_LC_7_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__16651\,
            in1 => \N__16604\,
            in2 => \_gnd_net_\,
            in3 => \N__16564\,
            lcout => \uu2.N_158\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.segmentUQ_0_5_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010100000110010"
        )
    port map (
            in0 => \N__19358\,
            in1 => \N__19311\,
            in2 => \N__19741\,
            in3 => \N__19269\,
            lcout => OPEN,
            ltout => \Lab_UT.segmentUQ_0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_90_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19886\,
            in2 => \N__16552\,
            in3 => \N__19559\,
            lcout => \uu2.bitmapZ0Z_90\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_90C_net\,
            ce => 'H',
            sr => \N__26045\
        );

    \Lab_UT.bcd2segment1.segment_1_6_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111100"
        )
    port map (
            in0 => \N__19357\,
            in1 => \N__19310\,
            in2 => \N__19740\,
            in3 => \N__19268\,
            lcout => \Lab_UT.segment_1_2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.segmentUQ_i_a4_1_6_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__19267\,
            in1 => \N__19737\,
            in2 => \N__19317\,
            in3 => \N__19360\,
            lcout => OPEN,
            ltout => \Lab_UT.N_65_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_186_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111011001100"
        )
    port map (
            in0 => \N__19560\,
            in1 => \N__19855\,
            in2 => \N__16825\,
            in3 => \N__16822\,
            lcout => \uu2.bitmapZ0Z_186\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_90C_net\,
            ce => 'H',
            sr => \N__26045\
        );

    \Lab_UT.bcd2segment1.segmentUQ_i_a3_4_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100000010"
        )
    port map (
            in0 => \N__19270\,
            in1 => \N__19736\,
            in2 => \N__19318\,
            in3 => \N__19359\,
            lcout => OPEN,
            ltout => \Lab_UT.N_76_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_218_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110111001100"
        )
    port map (
            in0 => \N__19327\,
            in1 => \N__19856\,
            in2 => \N__16807\,
            in3 => \N__19564\,
            lcout => \uu2.bitmapZ0Z_218\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_90C_net\,
            ce => 'H',
            sr => \N__26045\
        );

    \uu2.bitmap_RNICFK91_90_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001111"
        )
    port map (
            in0 => \N__16804\,
            in1 => \N__19435\,
            in2 => \N__16798\,
            in3 => \N__16767\,
            lcout => \uu2.bitmap_pmux_25_bm_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment2.segment_1_6_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111100"
        )
    port map (
            in0 => \N__20041\,
            in1 => \N__19983\,
            in2 => \N__19948\,
            in3 => \N__20071\,
            lcout => \Lab_UT.segment_1_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment2.segmentUQ_i_a3_4_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100000100"
        )
    port map (
            in0 => \N__20072\,
            in1 => \N__19937\,
            in2 => \N__19992\,
            in3 => \N__20042\,
            lcout => OPEN,
            ltout => \Lab_UT.N_76_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_212_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001110"
        )
    port map (
            in0 => \N__20166\,
            in1 => \N__19878\,
            in2 => \N__16702\,
            in3 => \N__16906\,
            lcout => \uu2.bitmapZ0Z_212\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_212C_net\,
            ce => 'H',
            sr => \N__26043\
        );

    \Lab_UT.bcd2segment2.segmentUQ_i_a4_1_6_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__20073\,
            in1 => \N__19933\,
            in2 => \N__19991\,
            in3 => \N__20043\,
            lcout => OPEN,
            ltout => \Lab_UT.N_65_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_180_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111011001100"
        )
    port map (
            in0 => \N__20165\,
            in1 => \N__19877\,
            in2 => \N__16687\,
            in3 => \N__16684\,
            lcout => \uu2.bitmapZ0Z_180\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_212C_net\,
            ce => 'H',
            sr => \N__26043\
        );

    \Lab_UT.bcd2segment2.segmentUQ_i_a3_0_4_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19979\,
            in2 => \_gnd_net_\,
            in3 => \N__20040\,
            lcout => \Lab_UT.N_77_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_84_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__19876\,
            in1 => \N__20164\,
            in2 => \_gnd_net_\,
            in3 => \N__19903\,
            lcout => \uu2.bitmapZ0Z_84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_212C_net\,
            ce => 'H',
            sr => \N__26043\
        );

    \Lab_UT.didp.Mtens_alarm.q_RNIO8T96_3_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001101111"
        )
    port map (
            in0 => \N__16834\,
            in1 => \N__16979\,
            in2 => \N__17044\,
            in3 => \N__16857\,
            lcout => \Lab_UT.L3_segment4_0_i_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment4.segmentUQ_i_a4_1_6_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__16937\,
            in1 => \N__17039\,
            in2 => \N__16998\,
            in3 => \N__19588\,
            lcout => \Lab_UT.N_65\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Mtens_alarm.q_RNI7VK11_3_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26833\,
            in1 => \N__25533\,
            in2 => \_gnd_net_\,
            in3 => \N__19664\,
            lcout => \Lab_UT.Mten_at_3\,
            ltout => \Lab_UT.Mten_at_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment4.segment_1_3_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011011111"
        )
    port map (
            in0 => \N__16858\,
            in1 => \N__17038\,
            in2 => \N__16873\,
            in3 => \N__16833\,
            lcout => \Lab_UT.segment_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment4.segmentUQ_0_o2_5_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110100000000"
        )
    port map (
            in0 => \N__25852\,
            in1 => \N__19665\,
            in2 => \N__26890\,
            in3 => \N__16935\,
            lcout => \Lab_UT.N_69_0\,
            ltout => \Lab_UT.N_69_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment4.segmentUQ_i_a3_0_2_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__16983\,
            in1 => \_gnd_net_\,
            in2 => \N__16849\,
            in3 => \N__17037\,
            lcout => \Lab_UT.N_92\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment4.segmentUQ_0_o3_5_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19587\,
            in2 => \_gnd_net_\,
            in3 => \N__16934\,
            lcout => \Lab_UT.N_67_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment4.segmentUQ_i_a3_2_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000000000000"
        )
    port map (
            in0 => \N__16936\,
            in1 => \N__17033\,
            in2 => \N__16999\,
            in3 => \N__19589\,
            lcout => \Lab_UT.N_91\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment4.segmentUQ_i_a4_3_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000100010"
        )
    port map (
            in0 => \N__17032\,
            in1 => \N__19590\,
            in2 => \_gnd_net_\,
            in3 => \N__16938\,
            lcout => \Lab_UT.N_83\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Mtens_alarm.q_RNI1PK11_0_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30038\,
            in1 => \N__25061\,
            in2 => \_gnd_net_\,
            in3 => \N__19645\,
            lcout => \Lab_UT.Mten_at_0\,
            ltout => \Lab_UT.Mten_at_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment4.segmentUQ_i_a3_0_4_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__16987\,
            in1 => \_gnd_net_\,
            in2 => \N__16951\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.N_77\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Mtens_alarm.q_RNI3RK11_1_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__27948\,
            in1 => \N__26354\,
            in2 => \_gnd_net_\,
            in3 => \N__19644\,
            lcout => \Lab_UT.Mten_at_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Mtens_alarm.q_0_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__25062\,
            in1 => \N__23014\,
            in2 => \_gnd_net_\,
            in3 => \N__29102\,
            lcout => \Lab_UT.di_AMtens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29401\,
            ce => 'H',
            sr => \N__26065\
        );

    \Lab_UT.didp.Mtens_alarm.q_1_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__28821\,
            in1 => \_gnd_net_\,
            in2 => \N__23020\,
            in3 => \N__26355\,
            lcout => \Lab_UT.di_AMtens_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29401\,
            ce => 'H',
            sr => \N__26065\
        );

    \Lab_UT.dictrl.currState_2_2_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__17725\,
            in1 => \N__17419\,
            in2 => \N__17083\,
            in3 => \N__17401\,
            lcout => \Lab_UT.dictrl.currStateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29401\,
            ce => 'H',
            sr => \N__26065\
        );

    \Lab_UT.dictrl.currState_0_ret_14_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21520\,
            in1 => \N__20653\,
            in2 => \N__20815\,
            in3 => \N__21034\,
            lcout => \Lab_UT.dictrl.un2_dicAlarmTrig\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29395\,
            ce => 'H',
            sr => \N__26067\
        );

    \Lab_UT.dictrl.currState_0_ret_3_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__21033\,
            in1 => \N__21521\,
            in2 => \N__20794\,
            in3 => \N__20634\,
            lcout => \Lab_UT.dictrl.r_Sone_init5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29395\,
            ce => 'H',
            sr => \N__26067\
        );

    \Lab_UT.dictrl.currState_0_ret_29_RNO_0_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101011101011"
        )
    port map (
            in0 => \N__21519\,
            in1 => \N__21032\,
            in2 => \N__20659\,
            in3 => \N__20747\,
            lcout => \Lab_UT.dictrl.g0_13_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_RNII4T093_0_2_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110011001101"
        )
    port map (
            in0 => \N__21028\,
            in1 => \N__21515\,
            in2 => \N__20792\,
            in3 => \N__20623\,
            lcout => \Lab_UT.dictrl.g0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_RNO_10_1_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101000001010"
        )
    port map (
            in0 => \N__21516\,
            in1 => \N__21030\,
            in2 => \N__20657\,
            in3 => \N__20742\,
            lcout => \Lab_UT.dictrl.g0_i_o4_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_RNII4T093_1_2_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__21029\,
            in1 => \N__21517\,
            in2 => \N__20793\,
            in3 => \N__20627\,
            lcout => \Lab_UT.dictrl.r_dicLdMtens16_reti\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_RNII4T093_2_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101110101011"
        )
    port map (
            in0 => \N__21518\,
            in1 => \N__21031\,
            in2 => \N__20658\,
            in3 => \N__20746\,
            lcout => \Lab_UT.dictrl.currState_0_ret_20and_1_0\,
            ltout => \Lab_UT.dictrl.currState_0_ret_20and_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_RNI82L3I6_2_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__24689\,
            in1 => \_gnd_net_\,
            in2 => \N__17116\,
            in3 => \N__20118\,
            lcout => \Lab_UT.dictrl.N_258_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.dicLdASones_RNI1C3E5_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__17364\,
            in1 => \N__20506\,
            in2 => \_gnd_net_\,
            in3 => \N__17374\,
            lcout => \Lab_UT.ld_enable_ASones\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_3_3_rep1_RNI2J197_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010100000"
        )
    port map (
            in0 => \N__17113\,
            in1 => \N__27802\,
            in2 => \N__20396\,
            in3 => \N__27544\,
            lcout => \Lab_UT.dictrl.N_13\,
            ltout => \Lab_UT.dictrl.N_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_3_3_rep1_RNIKKEKM_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__17724\,
            in1 => \N__17415\,
            in2 => \N__17404\,
            in3 => \N__17394\,
            lcout => \Lab_UT.dictrl.nextStateZ0Z_2\,
            ltout => \Lab_UT.dictrl.nextStateZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_3_3_rep1_RNI39J171_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001010"
        )
    port map (
            in0 => \N__21514\,
            in1 => \_gnd_net_\,
            in2 => \N__17377\,
            in3 => \N__24679\,
            lcout => \Lab_UT.dictrl.currState_ret_1and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_RNIMNQP4_2_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__27545\,
            in1 => \_gnd_net_\,
            in2 => \N__27814\,
            in3 => \N__23670\,
            lcout => \Lab_UT.dictrl.dicLdASones_rst\,
            ltout => \Lab_UT.dictrl.dicLdASones_rst_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.dicLdASones_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011100010"
        )
    port map (
            in0 => \N__17365\,
            in1 => \N__20507\,
            in2 => \N__17368\,
            in3 => \N__20560\,
            lcout => \Lab_UT.dictrl.dicLdASonesZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29391\,
            ce => 'H',
            sr => \N__23671\
        );

    \Lab_UT.dictrl.currState_2_RNIFK4DG_1_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24676\,
            in2 => \_gnd_net_\,
            in3 => \N__21513\,
            lcout => \Lab_UT.dictrl.N_5ctr\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_0_ret_1_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010001000000010"
        )
    port map (
            in0 => \N__21040\,
            in1 => \N__17308\,
            in2 => \N__17185\,
            in3 => \N__17266\,
            lcout => \Lab_UT.dictrl.r_Sone_init5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29385\,
            ce => 'H',
            sr => \N__26070\
        );

    \Lab_UT.dictrl.currState_0_ret_5_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000111010"
        )
    port map (
            in0 => \N__17307\,
            in1 => \N__17265\,
            in2 => \N__17183\,
            in3 => \N__21041\,
            lcout => \Lab_UT.dictrl.r_dicLdMtens14_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29385\,
            ce => 'H',
            sr => \N__26070\
        );

    \Lab_UT.dictrl.currState_2_RNIRPGDN_1_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011101111"
        )
    port map (
            in0 => \N__17264\,
            in1 => \N__24684\,
            in2 => \N__17184\,
            in3 => \N__17306\,
            lcout => \Lab_UT.dictrl.N_7ctr\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_RNI4F3LS1_1_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101000000000"
        )
    port map (
            in0 => \N__17305\,
            in1 => \N__17263\,
            in2 => \N__17182\,
            in3 => \N__21038\,
            lcout => \Lab_UT.dictrl.r_dicLdMtens15_1i\,
            ltout => \Lab_UT.dictrl.r_dicLdMtens15_1i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_RNI7OMM33_1_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__21574\,
            in1 => \N__24685\,
            in2 => \N__17602\,
            in3 => \N__20757\,
            lcout => \Lab_UT.dictrl.currState_ret_3and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_0_ret_28_RNO_3_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__20756\,
            in1 => \N__21573\,
            in2 => \_gnd_net_\,
            in3 => \N__21039\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.currState_0_ret_28_RNOZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_0_ret_28_RNO_1_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011110101111"
        )
    port map (
            in0 => \N__17587\,
            in1 => \N__17571\,
            in2 => \N__17491\,
            in3 => \N__17479\,
            lcout => \Lab_UT.dictrl.N_8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_RNIS2IML1_2_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__24683\,
            in1 => \N__21572\,
            in2 => \_gnd_net_\,
            in3 => \N__21037\,
            lcout => \Lab_UT.dictrl.r_dicLdMtens21_1_reti\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.decoder.g0_10_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__17710\,
            in1 => \N__17472\,
            in2 => \N__18186\,
            in3 => \N__17660\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.de_littleA_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__g0_3_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000001010"
        )
    port map (
            in0 => \N__20891\,
            in1 => \N__24217\,
            in2 => \N__17458\,
            in3 => \N__27748\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_37_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_RNIQ4BA8_1_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__17926\,
            in1 => \N__18070\,
            in2 => \N__17455\,
            in3 => \N__18055\,
            lcout => \Lab_UT.dictrl.g0_15_rn_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_3_3_rep1_RNIRM2Q_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__20394\,
            in1 => \N__25025\,
            in2 => \N__23458\,
            in3 => \N__17925\,
            lcout => \Lab_UT.dictrl.G_19_0_a7_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_2_rep1_es_RNIELCR_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__21703\,
            in1 => \N__21937\,
            in2 => \N__21780\,
            in3 => \N__17697\,
            lcout => \G_19_0_a7_4_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_RNIEPCJ_1_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18053\,
            in2 => \_gnd_net_\,
            in3 => \N__17924\,
            lcout => \Lab_UT.dictrl.currState_2_RNIEPCJZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_RNI2SKC_3_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__18088\,
            in1 => \N__23448\,
            in2 => \_gnd_net_\,
            in3 => \N__20393\,
            lcout => \Lab_UT.dictrl.N_1612_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_RNIEGFT_0_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__23452\,
            in1 => \N__18054\,
            in2 => \N__21268\,
            in3 => \N__17927\,
            lcout => \Lab_UT.dictrl.G_19_0_a7_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.decoder.g0_2_2_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__21832\,
            in1 => \N__21918\,
            in2 => \N__21991\,
            in3 => \N__17695\,
            lcout => \Lab_UT.dictrl.decoder.g0_2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.decoder.de_cr_2_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21891\,
            in2 => \_gnd_net_\,
            in3 => \N__17616\,
            lcout => \Lab_UT_dictrl_decoder_de_cr_2\,
            ltout => \Lab_UT_dictrl_decoder_de_cr_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.decoder.g0_4_3_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__21833\,
            in1 => \_gnd_net_\,
            in2 => \N__17701\,
            in3 => \N__17696\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.decoder.g0_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.decoder.g0_11_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21358\,
            in1 => \N__18172\,
            in2 => \N__17671\,
            in3 => \N__17667\,
            lcout => \Lab_UT.dictrl.de_cr_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_fast_2_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28906\,
            lcout => bu_rx_data_fast_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29377\,
            ce => \N__25423\,
            sr => \N__26097\
        );

    \buart.Z_rx.shifter_fast_1_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__28573\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_fast_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29377\,
            ce => \N__25423\,
            sr => \N__26097\
        );

    \Lab_UT.dictrl.decoder.g0_13_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18175\,
            in1 => \N__18409\,
            in2 => \N__18331\,
            in3 => \N__18367\,
            lcout => \Lab_UT.dictrl.de_cr_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.decoder.de_cr_1_1_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__24441\,
            in1 => \N__25300\,
            in2 => \N__24294\,
            in3 => \N__21414\,
            lcout => \Lab_UT_dictrl_decoder_de_cr_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.decoder.g0_17_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__25374\,
            in1 => \N__18307\,
            in2 => \N__29048\,
            in3 => \N__18273\,
            lcout => \Lab_UT.dictrl.decoder.g0_4Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.decoder.g0_16_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__28597\,
            in1 => \N__28924\,
            in2 => \_gnd_net_\,
            in3 => \N__18226\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.decoder.g0_3_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.decoder.g0_15_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18174\,
            in1 => \N__18385\,
            in2 => \N__18379\,
            in3 => \N__18366\,
            lcout => \Lab_UT.dictrl.de_cr_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.decoder.g0_14_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__18274\,
            in1 => \N__25375\,
            in2 => \N__18320\,
            in3 => \N__29026\,
            lcout => \Lab_UT.dictrl.decoder.g0_4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__g0_15_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__25373\,
            in1 => \N__18306\,
            in2 => \N__29047\,
            in3 => \N__18272\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__g0_12_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__24442\,
            in1 => \N__18225\,
            in2 => \N__18190\,
            in3 => \N__18173\,
            lcout => \Lab_UT.dictrl.g0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.uu0.l_count_6_LC_8_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001010101000000"
        )
    port map (
            in0 => \N__23233\,
            in1 => \N__22194\,
            in2 => \N__18517\,
            in3 => \N__22036\,
            lcout => \Lab_UT.uu0.l_countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29471\,
            ce => \N__22173\,
            sr => \N__26102\
        );

    \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_8_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__22035\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18513\,
            lcout => OPEN,
            ltout => \Lab_UT.uu0.un99_ci_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.uu0.l_count_7_LC_8_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001010101000000"
        )
    port map (
            in0 => \N__23234\,
            in1 => \N__22195\,
            in2 => \N__18520\,
            in3 => \N__18502\,
            lcout => \Lab_UT.uu0.l_countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29471\,
            ce => \N__22173\,
            sr => \N__26102\
        );

    \Lab_UT.uu0.l_count_16_LC_8_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__18621\,
            in1 => \N__22578\,
            in2 => \N__18609\,
            in3 => \N__23232\,
            lcout => \Lab_UT.uu0.l_countZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29471\,
            ce => \N__22173\,
            sr => \N__26102\
        );

    \Lab_UT.uu0.l_count_17_LC_8_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__22579\,
            in1 => \N__18601\,
            in2 => \N__18486\,
            in3 => \N__18622\,
            lcout => \Lab_UT.uu0.l_countZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29471\,
            ce => \N__22173\,
            sr => \N__26102\
        );

    \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_8_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22214\,
            in2 => \_gnd_net_\,
            in3 => \N__22128\,
            lcout => \Lab_UT.uu0.un88_ci_3\,
            ltout => \Lab_UT.uu0.un88_ci_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_8_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22192\,
            in1 => \N__22034\,
            in2 => \N__18505\,
            in3 => \N__18501\,
            lcout => \Lab_UT.uu0.un110_ci\,
            ltout => \Lab_UT.uu0.un110_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_8_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18620\,
            in1 => \N__18479\,
            in2 => \N__18463\,
            in3 => \N__22577\,
            lcout => \Lab_UT.uu0.un220_ci\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.uu0.l_count_10_LC_8_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__18555\,
            in1 => \N__18454\,
            in2 => \N__18608\,
            in3 => \N__18428\,
            lcout => \Lab_UT.uu0.l_countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29464\,
            ce => \N__22170\,
            sr => \N__26100\
        );

    \Lab_UT.uu0.l_count_RNIKE6P_2_LC_8_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__18427\,
            in1 => \N__18554\,
            in2 => \N__18671\,
            in3 => \N__22235\,
            lcout => OPEN,
            ltout => \Lab_UT.uu0.un4_l_count_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.uu0.l_count_RNIAK6Q1_4_LC_8_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__25200\,
            in1 => \N__22213\,
            in2 => \N__18700\,
            in3 => \N__18643\,
            lcout => \Lab_UT.uu0.un4_l_count_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.uu0.l_count_14_LC_8_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__18690\,
            in1 => \N__18646\,
            in2 => \N__18672\,
            in3 => \N__18593\,
            lcout => \Lab_UT.uu0.l_countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29464\,
            ce => \N__22170\,
            sr => \N__26100\
        );

    \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_8_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__18670\,
            in1 => \N__18689\,
            in2 => \_gnd_net_\,
            in3 => \N__18645\,
            lcout => OPEN,
            ltout => \Lab_UT.uu0.un187_ci_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.uu0.l_count_15_LC_8_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__22057\,
            in1 => \N__18594\,
            in2 => \N__18697\,
            in3 => \N__23223\,
            lcout => \Lab_UT.uu0.l_countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29464\,
            ce => \N__22170\,
            sr => \N__26100\
        );

    \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_8_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22056\,
            in1 => \N__18688\,
            in2 => \N__18673\,
            in3 => \N__18644\,
            lcout => \Lab_UT.uu0.un198_ci_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.uu0.l_count_8_LC_8_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18592\,
            in2 => \_gnd_net_\,
            in3 => \N__18556\,
            lcout => \Lab_UT.uu0.l_countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29464\,
            ce => \N__22170\,
            sr => \N__26100\
        );

    \uu2.w_addr_user_RNI0FES5_2_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22312\,
            in2 => \_gnd_net_\,
            in3 => \N__22423\,
            lcout => \uu2.un28_w_addr_user_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un1_w_user_lf_LC_8_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__18823\,
            in1 => \N__22280\,
            in2 => \N__25687\,
            in3 => \N__22827\,
            lcout => \uu2.un1_w_user_lf_0\,
            ltout => \uu2.un1_w_user_lf_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_RNIMJ3O2_2_LC_8_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__18891\,
            in1 => \N__26143\,
            in2 => \N__18523\,
            in3 => \N__18879\,
            lcout => \uu2.w_addr_user_RNIMJ3O2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vram_wr_en_0_i_LC_8_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100110011"
        )
    port map (
            in0 => \N__18880\,
            in1 => \N__29490\,
            in2 => \_gnd_net_\,
            in3 => \N__22294\,
            lcout => \uu2.vram_wr_en_0_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_RNIARA43_2_LC_8_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22293\,
            in1 => \N__18898\,
            in2 => \N__18892\,
            in3 => \N__18878\,
            lcout => \uu2.un28_w_addr_user_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un1_w_user_cr_LC_8_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__25683\,
            in1 => \N__18829\,
            in2 => \N__25594\,
            in3 => \N__22661\,
            lcout => \uu2.un1_w_user_cr_0\,
            ltout => \uu2.un1_w_user_cr_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un4_w_user_data_rdy_0_LC_8_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__22292\,
            in1 => \_gnd_net_\,
            in2 => \N__18868\,
            in3 => \_gnd_net_\,
            lcout => \uu2.un4_w_user_data_rdyZ0Z_0\,
            ltout => \uu2.un4_w_user_data_rdyZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_14_LC_8_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18863\,
            in2 => \N__18847\,
            in3 => \N__22281\,
            lcout => \uu2.mem0.w_data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un1_w_user_cr_4_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__22613\,
            in1 => \N__22632\,
            in2 => \N__22282\,
            in3 => \N__22820\,
            lcout => \uu2.un1_w_user_crZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un1_w_user_lf_4_LC_8_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__22631\,
            in1 => \N__25586\,
            in2 => \N__22665\,
            in3 => \N__22614\,
            lcout => \uu2.un1_w_user_lfZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_10_LC_8_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__18751\,
            in1 => \N__25590\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uu2.mem0.w_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__19062\,
            in1 => \N__18750\,
            in2 => \_gnd_net_\,
            in3 => \N__19495\,
            lcout => \uu2.mem0.w_addr_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_0_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19064\,
            in2 => \_gnd_net_\,
            in3 => \N__22424\,
            lcout => \uu2.w_addr_userZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_0C_net\,
            ce => 'H',
            sr => \N__22327\
        );

    \uu2.w_addr_user_1_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__22425\,
            in1 => \_gnd_net_\,
            in2 => \N__19069\,
            in3 => \N__18968\,
            lcout => \uu2.w_addr_userZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_0C_net\,
            ce => 'H',
            sr => \N__22327\
        );

    \uu2.w_addr_user_2_LC_8_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__18969\,
            in1 => \N__19068\,
            in2 => \N__19034\,
            in3 => \N__22426\,
            lcout => \uu2.w_addr_userZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_0C_net\,
            ce => 'H',
            sr => \N__22327\
        );

    \uu2.vbuf_w_addr_user.counter_gen_label_4__un404_ci_LC_8_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__19063\,
            in1 => \N__19023\,
            in2 => \N__18997\,
            in3 => \N__18967\,
            lcout => \uu2.un404_ci\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.curr_LED_1_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010101000000"
        )
    port map (
            in0 => \N__26151\,
            in1 => \N__29725\,
            in2 => \N__25456\,
            in3 => \N__29612\,
            lcout => \Lab_UT.didp.curr_LEDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29441\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.curr_LED_0_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__29724\,
            in1 => \N__25452\,
            in2 => \_gnd_net_\,
            in3 => \N__26152\,
            lcout => \Lab_UT.didp.curr_LEDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29441\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.uu0.counter_gen_label_3__un252_ci_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__19227\,
            in1 => \N__19239\,
            in2 => \_gnd_net_\,
            in3 => \N__19139\,
            lcout => OPEN,
            ltout => \resetGen.un252_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_3_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010100010000"
        )
    port map (
            in0 => \N__20424\,
            in1 => \N__19187\,
            in2 => \N__18940\,
            in3 => \N__18933\,
            lcout => \resetGen.reset_countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29441\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_1_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011000110"
        )
    port map (
            in0 => \N__19228\,
            in1 => \N__19240\,
            in2 => \N__19192\,
            in3 => \N__20422\,
            lcout => \resetGen.reset_countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29441\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.uu0.counter_gen_label_2__un241_ci_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__19238\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19226\,
            lcout => \resetGen.un241_ci\,
            ltout => \resetGen.un241_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_2_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010011100"
        )
    port map (
            in0 => \N__19186\,
            in1 => \N__19140\,
            in2 => \N__19147\,
            in3 => \N__20423\,
            lcout => \resetGen.reset_countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29441\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.uu0.delay_line_RNII8EF5_1_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__19123\,
            in1 => \N__22146\,
            in2 => \_gnd_net_\,
            in3 => \N__23235\,
            lcout => \Lab_UT.uu0.un11_l_count_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_93_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011110000"
        )
    port map (
            in0 => \N__19563\,
            in1 => \_gnd_net_\,
            in2 => \N__19887\,
            in3 => \N__19075\,
            lcout => \uu2.bitmapZ0Z_93\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_93C_net\,
            ce => 'H',
            sr => \N__26048\
        );

    \Lab_UT.didp.Sones_alarm.q_RNIOCVC5_1_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111010110101"
        )
    port map (
            in0 => \N__19354\,
            in1 => \N__19304\,
            in2 => \N__19738\,
            in3 => \N__19265\,
            lcout => \Lab_UT.L3_segment1_1_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Sones_alarm.q_RNIOCVC5_1_1_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000010000110"
        )
    port map (
            in0 => \N__19264\,
            in1 => \N__19355\,
            in2 => \N__19316\,
            in3 => \N__19726\,
            lcout => OPEN,
            ltout => \Lab_UT.L3_segment1_0_i_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_58_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19851\,
            in2 => \N__19087\,
            in3 => \N__19562\,
            lcout => \uu2.bitmapZ0Z_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_93C_net\,
            ce => 'H',
            sr => \N__26048\
        );

    \Lab_UT.didp.Sones_alarm.q_RNIOCVC5_2_1_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110111010111"
        )
    port map (
            in0 => \N__19263\,
            in1 => \N__19353\,
            in2 => \N__19315\,
            in3 => \N__19722\,
            lcout => \Lab_UT.L3_segment1_0_i_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Sones_alarm.q_RNIOCVC5_0_1_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101111101111"
        )
    port map (
            in0 => \N__19356\,
            in1 => \N__19305\,
            in2 => \N__19739\,
            in3 => \N__19266\,
            lcout => OPEN,
            ltout => \Lab_UT.L3_segment1_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_221_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__19561\,
            in1 => \_gnd_net_\,
            in2 => \N__19522\,
            in3 => \N__19857\,
            lcout => \uu2.bitmapZ0Z_221\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_93C_net\,
            ce => 'H',
            sr => \N__26048\
        );

    \uu2.bitmap_RNI1D952_93_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000110011"
        )
    port map (
            in0 => \N__19519\,
            in1 => \N__19513\,
            in2 => \N__19507\,
            in3 => \N__19491\,
            lcout => \uu2.bitmap_RNI1D952Z0Z_93\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.dicLdAStens_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__20515\,
            in1 => \N__20457\,
            in2 => \N__20476\,
            in3 => \N__20569\,
            lcout => \Lab_UT.dictrl.dicLdAStensZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29426\,
            ce => 'H',
            sr => \N__23899\
        );

    \Lab_UT.didp.Sones_alarm.q_RNI3O7B1_0_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29820\,
            in1 => \N__23075\,
            in2 => \_gnd_net_\,
            in3 => \N__19666\,
            lcout => \Lab_UT.Sone_at_0\,
            ltout => \Lab_UT.Sone_at_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.segmentUQ_i_a3_0_4_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19330\,
            in3 => \N__19306\,
            lcout => \Lab_UT.N_77_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Sones_alarm.q_RNI9U7B1_3_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26188\,
            in1 => \N__22925\,
            in2 => \_gnd_net_\,
            in3 => \N__19669\,
            lcout => \Lab_UT.Sone_at_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Sones_alarm.q_RNI7S7B1_2_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__19667\,
            in1 => \N__26229\,
            in2 => \_gnd_net_\,
            in3 => \N__23036\,
            lcout => \Lab_UT.Sone_at_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Stens_alarm.q_RNIHF5B1_2_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25625\,
            in1 => \N__27162\,
            in2 => \_gnd_net_\,
            in3 => \N__19670\,
            lcout => \Lab_UT.Sten_at_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Stens_alarm.q_RNIDB5B1_0_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__19668\,
            in1 => \N__29689\,
            in2 => \_gnd_net_\,
            in3 => \N__25724\,
            lcout => \Lab_UT.Sten_at_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Stens_alarm.q_RNIJH5B1_3_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__27126\,
            in1 => \N__22979\,
            in2 => \_gnd_net_\,
            in3 => \N__19671\,
            lcout => \Lab_UT.Sten_at_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Stens_alarm.q_RNIFD5B1_1_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__19660\,
            in1 => \_gnd_net_\,
            in2 => \N__25809\,
            in3 => \N__27872\,
            lcout => \Lab_UT.Sten_at_1\,
            ltout => \Lab_UT.Sten_at_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment2.segmentUQ_0_5_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010100000110010"
        )
    port map (
            in0 => \N__20030\,
            in1 => \N__19987\,
            in2 => \N__19954\,
            in3 => \N__19923\,
            lcout => \Lab_UT.segmentUQ_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_0_ret_11_RNIA2D93_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__20824\,
            in1 => \N__27811\,
            in2 => \_gnd_net_\,
            in3 => \N__27300\,
            lcout => \Lab_UT.dicLdStens_latmux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_0_ret_14_RNID3D61_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__26675\,
            in1 => \N__24172\,
            in2 => \N__29491\,
            in3 => \N__23646\,
            lcout => \Lab_UT.dictrl.L3_segment1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Sones_alarm.q_RNI5Q7B1_1_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__23059\,
            in1 => \N__28104\,
            in2 => \_gnd_net_\,
            in3 => \N__19659\,
            lcout => \Lab_UT.Sone_at_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_0_ret_3_RNI9MVL_0_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__26676\,
            in1 => \N__23476\,
            in2 => \_gnd_net_\,
            in3 => \N__23161\,
            lcout => \Lab_UT.dictrl.r_enable1_2_i_m\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.r_alarm_or_time_RNI9J3I_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__24157\,
            in1 => \N__23637\,
            in2 => \_gnd_net_\,
            in3 => \N__20223\,
            lcout => \Lab_UT.alarm_or_time_0\,
            ltout => \Lab_UT.alarm_or_time_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Mtens_alarm.q_RNI5TK11_2_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__25844\,
            in1 => \_gnd_net_\,
            in2 => \N__19612\,
            in3 => \N__26873\,
            lcout => \Lab_UT.Mten_at_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.dicLdStens_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011110000"
        )
    port map (
            in0 => \N__29939\,
            in1 => \N__23092\,
            in2 => \N__23113\,
            in3 => \N__29882\,
            lcout => \Lab_UT.dicLdStens\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29409\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_0_ret_3_RNI9MVL_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__26677\,
            in1 => \N__23477\,
            in2 => \_gnd_net_\,
            in3 => \N__23162\,
            lcout => \Lab_UT.dictrl.r_enable1_2_m\,
            ltout => \Lab_UT.dictrl.r_enable1_2_m_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.r_enable2_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101010001"
        )
    port map (
            in0 => \N__23440\,
            in1 => \N__20260\,
            in2 => \N__20191\,
            in3 => \N__20179\,
            lcout => \Lab_UT.dictrl.r_enableZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29409\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_0_ret_29_RNIPGJ2_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23439\,
            in2 => \_gnd_net_\,
            in3 => \N__26149\,
            lcout => \Lab_UT.dictrl.g0_i_a4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.r_enable2_RNI8DR61_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__24158\,
            in1 => \N__20178\,
            in2 => \N__23170\,
            in3 => \N__23638\,
            lcout => \Lab_UT.dictrl.enableSeg2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_0_ret_22_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__20125\,
            in1 => \N__24687\,
            in2 => \_gnd_net_\,
            in3 => \N__20119\,
            lcout => \Lab_UT.un1_r_Sone_init5_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29402\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_ret_0_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__24686\,
            in1 => \N__20767\,
            in2 => \N__24730\,
            in3 => \N__21606\,
            lcout => \Lab_UT.dictrl.r_dicLdMtens19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29402\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_0_ret_23_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__20561\,
            in1 => \N__24726\,
            in2 => \_gnd_net_\,
            in3 => \N__24688\,
            lcout => \Lab_UT.dictrl.r_dicLdMtens23_i_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29402\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.r_enable2_RNO_1_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__20086\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20206\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.r_enable2_3_iv_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.r_enable2_RNO_0_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20212\,
            in1 => \N__20235\,
            in2 => \N__20263\,
            in3 => \N__23595\,
            lcout => \Lab_UT.dictrl.r_enable2_3_iv_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.r_alarm_or_time_RNO_0_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20251\,
            in2 => \_gnd_net_\,
            in3 => \N__20236\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.un1_r_dicLdMtens19_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.r_alarm_or_time_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010100000001"
        )
    port map (
            in0 => \N__23478\,
            in1 => \N__23435\,
            in2 => \N__20227\,
            in3 => \N__20224\,
            lcout => \Lab_UT.dictrl.r_alarm_or_timeZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29402\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_0_ret_12_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__21615\,
            in1 => \N__20661\,
            in2 => \N__20806\,
            in3 => \N__21095\,
            lcout => \Lab_UT.dictrl.r_dicLdMtens15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29396\,
            ce => 'H',
            sr => \N__26071\
        );

    \Lab_UT.dictrl.currState_0_ret_16_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__21091\,
            in1 => \N__21619\,
            in2 => \N__20810\,
            in3 => \N__20665\,
            lcout => \Lab_UT.dictrl.r_dicLdMtens18_i_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29396\,
            ce => 'H',
            sr => \N__26071\
        );

    \Lab_UT.dictrl.currState_0_ret_18_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__21616\,
            in1 => \N__20662\,
            in2 => \N__20807\,
            in3 => \N__21096\,
            lcout => \Lab_UT.dictrl.r_dicLdMtens17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29396\,
            ce => 'H',
            sr => \N__26071\
        );

    \Lab_UT.dictrl.currState_0_ret_19_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__21092\,
            in1 => \N__21620\,
            in2 => \N__20811\,
            in3 => \N__20666\,
            lcout => \Lab_UT.dictrl.r_dicLdMtens17_i_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29396\,
            ce => 'H',
            sr => \N__26071\
        );

    \Lab_UT.dictrl.currState_0_ret_6_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__21617\,
            in1 => \N__20663\,
            in2 => \N__20808\,
            in3 => \N__21097\,
            lcout => \Lab_UT.dictrl.r_dicLdMtens14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29396\,
            ce => 'H',
            sr => \N__26071\
        );

    \Lab_UT.dictrl.currState_0_ret_7_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__21093\,
            in1 => \N__21621\,
            in2 => \N__20812\,
            in3 => \N__20667\,
            lcout => \Lab_UT.dictrl.r_dicLdMtens14_i_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29396\,
            ce => 'H',
            sr => \N__26071\
        );

    \Lab_UT.dictrl.currState_0_ret_11_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__21614\,
            in1 => \N__20660\,
            in2 => \N__20805\,
            in3 => \N__21094\,
            lcout => \Lab_UT.dictrl.r_dicLdMtens16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29396\,
            ce => 'H',
            sr => \N__26071\
        );

    \Lab_UT.dictrl.currState_0_ret_15_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__21090\,
            in1 => \N__21618\,
            in2 => \N__20809\,
            in3 => \N__20664\,
            lcout => \Lab_UT.dictrl.un2_dicAlarmTrig_i_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29396\,
            ce => 'H',
            sr => \N__26071\
        );

    \Lab_UT.dictrl.currState_0_ret_18_RNIH2D93_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__20578\,
            in1 => \N__27806\,
            in2 => \_gnd_net_\,
            in3 => \N__27559\,
            lcout => \Lab_UT.dicLdSones_latmux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.dicLdAMones_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__20562\,
            in1 => \N__20530\,
            in2 => \N__20539\,
            in3 => \N__20518\,
            lcout => \Lab_UT.dictrl.dicLdAMonesZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29392\,
            ce => 'H',
            sr => \N__23920\
        );

    \Lab_UT.dictrl.currState_ret_7_RNIUEJQ4_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__23913\,
            in1 => \N__27807\,
            in2 => \_gnd_net_\,
            in3 => \N__27560\,
            lcout => \Lab_UT.dictrl.dicLdAMones_rst\,
            ltout => \Lab_UT.dictrl.dicLdAMones_rst_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.dicLdAMones_RNI3BNL5_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20529\,
            in2 => \N__20521\,
            in3 => \N__20517\,
            lcout => \Lab_UT.ld_enable_AMones\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.dicLdAStens_RNI7OAH5_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__20516\,
            in1 => \N__20475\,
            in2 => \_gnd_net_\,
            in3 => \N__20458\,
            lcout => \Lab_UT.ld_enable_AStens\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.escKey_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__27808\,
            in1 => \N__21118\,
            in2 => \_gnd_net_\,
            in3 => \N__25435\,
            lcout => \resetGen.escKeyZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__m5_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101101010101"
        )
    port map (
            in0 => \N__20395\,
            in1 => \N__24476\,
            in2 => \_gnd_net_\,
            in3 => \N__20299\,
            lcout => \Lab_UT.dictrl.N_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.r_enable3_RNO_0_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__21325\,
            in1 => \N__21319\,
            in2 => \_gnd_net_\,
            in3 => \N__23686\,
            lcout => \Lab_UT.dictrl.r_enable3_3_iv_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_RNI86KI_6_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24295\,
            in2 => \_gnd_net_\,
            in3 => \N__28508\,
            lcout => OPEN,
            ltout => \buart.Z_rx.G_30_0_o3_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_RNIV4BN3_7_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__21634\,
            in1 => \N__25395\,
            in2 => \N__21295\,
            in3 => \N__21292\,
            lcout => OPEN,
            ltout => \N_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_0_ret_21_RNI88818_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000010001111"
        )
    port map (
            in0 => \N__21260\,
            in1 => \N__24475\,
            in2 => \N__21136\,
            in3 => \N__24011\,
            lcout => \Lab_UT.dictrl.N_21_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.escKey_4_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__28509\,
            in1 => \N__24447\,
            in2 => \N__24310\,
            in3 => \N__25396\,
            lcout => \resetGen.escKey_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_0_rep2_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24695\,
            in2 => \_gnd_net_\,
            in3 => \N__21107\,
            lcout => \Lab_UT.dictrl.currState_0_rep2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29386\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__g0_14_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__28743\,
            in1 => \N__28507\,
            in2 => \N__28947\,
            in3 => \N__25304\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__g0_7_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24296\,
            in1 => \N__20900\,
            in2 => \N__20860\,
            in3 => \N__24890\,
            lcout => \Lab_UT.dictrl.g0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.decoder.de_littleL_4_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21442\,
            in1 => \N__21346\,
            in2 => \N__21831\,
            in3 => \N__20838\,
            lcout => \Lab_UT.dictrl.de_littleL_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__g1_6_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__21347\,
            in1 => \N__21443\,
            in2 => \N__21781\,
            in3 => \N__21819\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g1_5_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__g1_2_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__21407\,
            in1 => \N__21649\,
            in2 => \N__21718\,
            in3 => \N__24308\,
            lcout => \Lab_UT.dictrl.g1_7_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_1_3_0__g1_3_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__21640\,
            in1 => \N__21699\,
            in2 => \_gnd_net_\,
            in3 => \N__21924\,
            lcout => \Lab_UT.dictrl.g1_4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_3_fast_3_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24704\,
            in2 => \_gnd_net_\,
            in3 => \N__21623\,
            lcout => \Lab_UT.dictrl.currState_fast_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29382\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_RNID9851_4_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__24443\,
            in1 => \N__28753\,
            in2 => \N__28964\,
            in3 => \N__25303\,
            lcout => \buart.Z_rx.G_30_0_o3_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_3_3_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24703\,
            in2 => \_gnd_net_\,
            in3 => \N__21622\,
            lcout => \Lab_UT.dictrl.currStateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29382\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.decoder.g0_12_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21445\,
            in1 => \N__21925\,
            in2 => \N__21987\,
            in3 => \N__21406\,
            lcout => \Lab_UT.dictrl.decoder.g0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_0_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28771\,
            lcout => bu_rx_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29378\,
            ce => \N__25424\,
            sr => \N__26101\
        );

    \buart.Z_rx.shifter_0_rep1_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28772\,
            lcout => bu_rx_data_0_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29378\,
            ce => \N__25424\,
            sr => \N__26101\
        );

    \buart.Z_rx.shifter_6_rep1_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25377\,
            lcout => bu_rx_data_6_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29378\,
            ce => \N__25424\,
            sr => \N__26101\
        );

    \buart.Z_rx.shifter_3_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25301\,
            lcout => bu_rx_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29378\,
            ce => \N__25424\,
            sr => \N__26101\
        );

    \buart.Z_rx.shifter_5_rep1_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24300\,
            lcout => bu_rx_data_5_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29378\,
            ce => \N__25424\,
            sr => \N__26101\
        );

    \buart.Z_rx.shifter_fast_3_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25302\,
            lcout => bu_rx_data_fast_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29378\,
            ce => \N__25424\,
            sr => \N__26101\
        );

    \buart.Z_rx.shifter_7_rep1_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21876\,
            lcout => bu_rx_data_7_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29378\,
            ce => \N__25424\,
            sr => \N__26101\
        );

    \Lab_UT.uu0.l_count_1_LC_9_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__22093\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22521\,
            lcout => \Lab_UT.uu0.l_countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29476\,
            ce => \N__22171\,
            sr => \N__26105\
        );

    \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_1_LC_9_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__22519\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22092\,
            lcout => \Lab_UT.uu0.un44_ci\,
            ltout => \Lab_UT.uu0.un44_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.uu0.l_count_3_LC_9_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__22243\,
            in1 => \N__22260\,
            in2 => \N__21784\,
            in3 => \N__23222\,
            lcout => \Lab_UT.uu0.l_countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29476\,
            ce => \N__22171\,
            sr => \N__26105\
        );

    \Lab_UT.uu0.l_count_0_LC_9_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22520\,
            in2 => \_gnd_net_\,
            in3 => \N__23220\,
            lcout => \Lab_UT.uu0.l_countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29476\,
            ce => \N__22171\,
            sr => \N__26105\
        );

    \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_9_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22259\,
            in1 => \N__22242\,
            in2 => \N__22522\,
            in3 => \N__22091\,
            lcout => \Lab_UT.uu0.un66_ci\,
            ltout => \Lab_UT.uu0.un66_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.uu0.l_count_4_LC_9_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22215\,
            in2 => \N__22219\,
            in3 => \N__23221\,
            lcout => \Lab_UT.uu0.l_countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29476\,
            ce => \N__22171\,
            sr => \N__26105\
        );

    \Lab_UT.uu0.l_count_5_LC_9_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__22216\,
            in1 => \N__22193\,
            in2 => \_gnd_net_\,
            in3 => \N__22129\,
            lcout => \Lab_UT.uu0.l_countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29476\,
            ce => \N__22171\,
            sr => \N__26105\
        );

    \Lab_UT.uu0.delay_line_0_LC_9_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22594\,
            in1 => \N__25210\,
            in2 => \N__22111\,
            in3 => \N__22537\,
            lcout => \Lab_UT.uu0.delay_lineZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29472\,
            ce => 'H',
            sr => \N__26104\
        );

    \Lab_UT.uu0.l_precount_3_LC_9_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__22539\,
            in1 => \N__22109\,
            in2 => \N__25216\,
            in3 => \N__22597\,
            lcout => \Lab_UT.uu0.l_precountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29472\,
            ce => 'H',
            sr => \N__26104\
        );

    \Lab_UT.uu0.l_count_RNIS3Q51_5_LC_9_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__22593\,
            in1 => \N__22127\,
            in2 => \N__22110\,
            in3 => \N__22090\,
            lcout => OPEN,
            ltout => \Lab_UT.uu0.un4_l_count_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.uu0.l_count_RNIC7FP1_18_LC_9_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22075\,
            in1 => \N__22055\,
            in2 => \N__22039\,
            in3 => \N__22033\,
            lcout => OPEN,
            ltout => \Lab_UT.uu0.un4_l_count_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.uu0.l_count_RNIRSCC5_3_LC_9_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22498\,
            in1 => \N__22018\,
            in2 => \N__22009\,
            in3 => \N__22006\,
            lcout => \Lab_UT.uu0.un4_l_count_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.uu0.l_precount_1_LC_9_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__25211\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22595\,
            lcout => \Lab_UT.uu0.l_precountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29472\,
            ce => 'H',
            sr => \N__26104\
        );

    \Lab_UT.uu0.l_precount_2_LC_9_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__22596\,
            in1 => \N__25212\,
            in2 => \_gnd_net_\,
            in3 => \N__22538\,
            lcout => \Lab_UT.uu0.l_precountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29472\,
            ce => 'H',
            sr => \N__26104\
        );

    \Lab_UT.uu0.l_count_RNIM5011_11_LC_9_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__22576\,
            in1 => \N__22556\,
            in2 => \N__22540\,
            in3 => \N__22515\,
            lcout => \Lab_UT.uu0.un4_l_count_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_5_LC_9_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__22428\,
            in1 => \N__22396\,
            in2 => \N__22462\,
            in3 => \N__22486\,
            lcout => \uu2.w_addr_userZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_5C_net\,
            ce => 'H',
            sr => \N__22326\
        );

    \uu2.w_addr_user_4_LC_9_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__22395\,
            in1 => \N__22455\,
            in2 => \_gnd_net_\,
            in3 => \N__22427\,
            lcout => \uu2.w_addr_userZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_5C_net\,
            ce => 'H',
            sr => \N__22326\
        );

    \uu2.w_addr_user_6_LC_9_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__22429\,
            in1 => \N__22397\,
            in2 => \N__22378\,
            in3 => \N__22350\,
            lcout => \uu2.w_addr_userZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_5C_net\,
            ce => 'H',
            sr => \N__22326\
        );

    \Lab_UT.display.cnt_RNIFA8M_0_2_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26511\,
            in2 => \_gnd_net_\,
            in3 => \N__26426\,
            lcout => \Lab_UT.display.N_150\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.display.rdy_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26428\,
            in1 => \N__26337\,
            in2 => \N__26515\,
            in3 => \N__26734\,
            lcout => \L3_tx_data_rdy\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29457\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.display.dOut_6_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__27424\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22854\,
            lcout => \L3_tx_data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29457\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.display.cnt_RNI5EC11_0_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25565\,
            in2 => \_gnd_net_\,
            in3 => \N__26335\,
            lcout => \Lab_UT.display.N_88\,
            ltout => \Lab_UT.display.N_88_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.display.dOut_1_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001110"
        )
    port map (
            in0 => \N__23131\,
            in1 => \N__25753\,
            in2 => \N__22669\,
            in3 => \N__22888\,
            lcout => \L3_tx_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29457\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.display.dOut_RNO_0_4_LC_9_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27367\,
            in2 => \_gnd_net_\,
            in3 => \N__25566\,
            lcout => OPEN,
            ltout => \Lab_UT.display.N_120_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.display.dOut_4_LC_9_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000011"
        )
    port map (
            in0 => \N__26336\,
            in1 => \N__25551\,
            in2 => \N__22642\,
            in3 => \N__26427\,
            lcout => \L3_tx_data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29457\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.display.dOut_5_LC_9_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010100010001"
        )
    port map (
            in0 => \N__25552\,
            in1 => \N__25567\,
            in2 => \N__26341\,
            in3 => \N__23614\,
            lcout => \L3_tx_data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29457\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.display.dOut_RNO_1_2_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110010"
        )
    port map (
            in0 => \N__26542\,
            in1 => \N__22733\,
            in2 => \N__22881\,
            in3 => \N__23037\,
            lcout => \Lab_UT.display.dOutP_0_iv_i_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.display.dOut_RNO_1_0_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011001110"
        )
    port map (
            in0 => \N__26541\,
            in1 => \N__22874\,
            in2 => \N__22764\,
            in3 => \N__23076\,
            lcout => \Lab_UT.display.dOutP_0_iv_i_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.display.cnt_RNIFA8M_1_2_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26509\,
            in2 => \_gnd_net_\,
            in3 => \N__26425\,
            lcout => \Lab_UT.display.N_153\,
            ltout => \Lab_UT.display.N_153_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.display.dOut_RNO_1_3_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011001100"
        )
    port map (
            in0 => \N__22984\,
            in1 => \N__25504\,
            in2 => \N__22600\,
            in3 => \N__26332\,
            lcout => \Lab_UT.display.dOutP_0_iv_i_2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.display.dOut_RNO_1_1_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011001100"
        )
    port map (
            in0 => \N__26331\,
            in1 => \N__26257\,
            in2 => \N__22882\,
            in3 => \N__23057\,
            lcout => \Lab_UT.display.dOutP_0_iv_i_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.display.dOut_RNO_2_3_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26333\,
            in2 => \_gnd_net_\,
            in3 => \N__22930\,
            lcout => OPEN,
            ltout => \Lab_UT.display.N_101_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.display.dOut_RNO_0_3_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__22873\,
            in1 => \N__26540\,
            in2 => \N__22861\,
            in3 => \N__22688\,
            lcout => OPEN,
            ltout => \Lab_UT.display.dOutP_0_iv_i_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.display.dOut_3_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001110"
        )
    port map (
            in0 => \N__23130\,
            in1 => \N__22858\,
            in2 => \N__22843\,
            in3 => \N__22840\,
            lcout => \L3_tx_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29450\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_addr_5_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__25108\,
            in1 => \N__25180\,
            in2 => \N__22792\,
            in3 => \N__25147\,
            lcout => \uu2.r_addrZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29442\,
            ce => 'H',
            sr => \N__26072\
        );

    \Lab_UT.didp.Mones_alarm.q_0_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__22711\,
            in1 => \N__22760\,
            in2 => \_gnd_net_\,
            in3 => \N__29103\,
            lcout => \Lab_UT.di_AMones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29442\,
            ce => 'H',
            sr => \N__26072\
        );

    \Lab_UT.didp.Mones_alarm.q_1_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28795\,
            in1 => \N__25775\,
            in2 => \_gnd_net_\,
            in3 => \N__22712\,
            lcout => \Lab_UT.di_AMones_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29442\,
            ce => 'H',
            sr => \N__26072\
        );

    \Lab_UT.didp.Mones_alarm.q_2_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__22713\,
            in1 => \N__22734\,
            in2 => \_gnd_net_\,
            in3 => \N__28610\,
            lcout => \Lab_UT.di_AMones_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29442\,
            ce => 'H',
            sr => \N__26072\
        );

    \Lab_UT.didp.Mones_alarm.q_3_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28983\,
            in1 => \N__22689\,
            in2 => \_gnd_net_\,
            in3 => \N__22714\,
            lcout => \Lab_UT.di_AMones_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29442\,
            ce => 'H',
            sr => \N__26072\
        );

    \Lab_UT.didp.Sones_alarm.q_0_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__22961\,
            in1 => \N__23077\,
            in2 => \_gnd_net_\,
            in3 => \N__29104\,
            lcout => \Lab_UT.di_ASones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29442\,
            ce => 'H',
            sr => \N__26072\
        );

    \Lab_UT.didp.Sones_alarm.q_1_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28796\,
            in1 => \N__23058\,
            in2 => \_gnd_net_\,
            in3 => \N__22962\,
            lcout => \Lab_UT.di_ASones_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29442\,
            ce => 'H',
            sr => \N__26072\
        );

    \Lab_UT.didp.Sones_alarm.q_2_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__22963\,
            in1 => \N__23038\,
            in2 => \_gnd_net_\,
            in3 => \N__28611\,
            lcout => \Lab_UT.di_ASones_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29442\,
            ce => 'H',
            sr => \N__26072\
        );

    \Lab_UT.didp.Mtens_alarm.q_2_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__23018\,
            in1 => \N__28608\,
            in2 => \_gnd_net_\,
            in3 => \N__25843\,
            lcout => \Lab_UT.di_AMtens_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29436\,
            ce => 'H',
            sr => \N__26069\
        );

    \Lab_UT.didp.Mtens_alarm.q_3_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__23019\,
            in1 => \N__25526\,
            in2 => \_gnd_net_\,
            in3 => \N__28985\,
            lcout => \Lab_UT.di_AMtens_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29436\,
            ce => 'H',
            sr => \N__26069\
        );

    \Lab_UT.didp.Stens_alarm.q_2_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25629\,
            in1 => \N__28609\,
            in2 => \_gnd_net_\,
            in3 => \N__22908\,
            lcout => \Lab_UT.di_AStens_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29436\,
            ce => 'H',
            sr => \N__26069\
        );

    \Lab_UT.didp.Stens_alarm.q_3_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__22909\,
            in1 => \N__22983\,
            in2 => \_gnd_net_\,
            in3 => \N__28986\,
            lcout => \Lab_UT.di_AStens_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29436\,
            ce => 'H',
            sr => \N__26069\
        );

    \Lab_UT.didp.Sones_alarm.q_3_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__28984\,
            in1 => \N__22953\,
            in2 => \_gnd_net_\,
            in3 => \N__22929\,
            lcout => \Lab_UT.di_ASones_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29436\,
            ce => 'H',
            sr => \N__26069\
        );

    \Lab_UT.didp.Stens_alarm.q_0_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__22906\,
            in1 => \N__25728\,
            in2 => \_gnd_net_\,
            in3 => \N__29105\,
            lcout => \Lab_UT.di_AStens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29436\,
            ce => 'H',
            sr => \N__26069\
        );

    \Lab_UT.didp.Stens_alarm.q_1_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28816\,
            in1 => \N__25802\,
            in2 => \_gnd_net_\,
            in3 => \N__22907\,
            lcout => \Lab_UT.di_AStens_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29436\,
            ce => 'H',
            sr => \N__26069\
        );

    \Lab_UT.uu0.sec_clk_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__23246\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23157\,
            lcout => \Lab_UT.halfPulse\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29436\,
            ce => 'H',
            sr => \N__26069\
        );

    \Lab_UT.didp.Stens_subtractor.q_7_i_o2_2_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110101111111"
        )
    port map (
            in0 => \N__28180\,
            in1 => \N__29959\,
            in2 => \N__23112\,
            in3 => \N__23091\,
            lcout => \Lab_UT.didp.Stens_subtractor.N_86\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.displayAlarm_1_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29540\,
            lcout => \Lab_UT.displayAlarmZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29427\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.dicLdStens_RNIQVHE3_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__23105\,
            in1 => \N__29958\,
            in2 => \_gnd_net_\,
            in3 => \N__23090\,
            lcout => \Lab_UT.ld_enable_Stens\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Stens_subtractor.q_RNI8PD76_1_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000010001"
        )
    port map (
            in0 => \N__26620\,
            in1 => \N__29683\,
            in2 => \_gnd_net_\,
            in3 => \N__27873\,
            lcout => \Lab_UT.didp.Stens_subtractor.q_RNI8PD76Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Stens_subtractor.q_RNIBBF11_2_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__26233\,
            in1 => \N__29761\,
            in2 => \_gnd_net_\,
            in3 => \N__27161\,
            lcout => \Lab_UT.didp.q_RNIBBF11_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Stens_subtractor.q_RNO_0_3_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110011001001"
        )
    port map (
            in0 => \N__26623\,
            in1 => \N__27118\,
            in2 => \N__26602\,
            in3 => \N__27159\,
            lcout => \Lab_UT.didp.Stens_subtractor.q_RNO_0_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Stens_subtractor.q_RNO_0_2_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000001"
        )
    port map (
            in0 => \N__29685\,
            in1 => \N__26622\,
            in2 => \N__27877\,
            in3 => \N__27160\,
            lcout => \Lab_UT.didp.Stens_subtractor.q_RNO_0_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Stens_subtractor.q_RNO_0_0_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100110011001"
        )
    port map (
            in0 => \N__26621\,
            in1 => \N__29684\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.didp.Stens_subtractor.un1_q_axb0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Stens_subtractor.q_0_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110101110101"
        )
    port map (
            in0 => \N__26969\,
            in1 => \N__23549\,
            in2 => \N__29106\,
            in3 => \N__23563\,
            lcout => \Lab_UT.didp.di_Stens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29417\,
            ce => 'H',
            sr => \N__28448\
        );

    \Lab_UT.didp.Stens_subtractor.q_3_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__23551\,
            in1 => \N__23557\,
            in2 => \N__28995\,
            in3 => \N__26971\,
            lcout => \Lab_UT.didp.di_Stens_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29417\,
            ce => 'H',
            sr => \N__28448\
        );

    \Lab_UT.didp.Stens_subtractor.q_2_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110101110101"
        )
    port map (
            in0 => \N__26970\,
            in1 => \N__23550\,
            in2 => \N__28612\,
            in3 => \N__23539\,
            lcout => \Lab_UT.didp.di_Stens_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29417\,
            ce => 'H',
            sr => \N__28448\
        );

    \Lab_UT.didp.Stens_subtractor.q_RNIDDF11_3_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__27119\,
            in1 => \_gnd_net_\,
            in2 => \N__29779\,
            in3 => \N__26197\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.q_RNIDDF11_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.curr_LED_RNIRNM52_1_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__29630\,
            in1 => \_gnd_net_\,
            in2 => \N__23533\,
            in3 => \N__23518\,
            lcout => led_c_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Mones_subtractor.q_RNI1TVP_3_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__26832\,
            in1 => \_gnd_net_\,
            in2 => \N__29778\,
            in3 => \N__28252\,
            lcout => \Lab_UT.didp.q_RNI1TVP_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.curr_LED_RNINJM52_1_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__23512\,
            in1 => \N__23506\,
            in2 => \_gnd_net_\,
            in3 => \N__29629\,
            lcout => led_c_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.r_dicRun_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000000101"
        )
    port map (
            in0 => \N__23482\,
            in1 => \N__26667\,
            in2 => \N__24742\,
            in3 => \N__23456\,
            lcout => \Lab_UT.ld_enable_dicRun\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29410\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_al_0_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__23572\,
            in1 => \N__23605\,
            in2 => \N__24121\,
            in3 => \N__26156\,
            lcout => \Lab_UT.dictrl.nextState_al_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29410\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.r_dicAlarmArmed_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000000110011"
        )
    port map (
            in0 => \N__29576\,
            in1 => \N__29126\,
            in2 => \N__27395\,
            in3 => \N__24058\,
            lcout => \Lab_UT.alarm_armed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29410\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.r_dicAlarmTrig_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000000010"
        )
    port map (
            in0 => \N__24057\,
            in1 => \N__29577\,
            in2 => \N__29130\,
            in3 => \N__23645\,
            lcout => \Lab_UT.dictrl.r_dicAlarmTrigZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29410\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.displayAlarm_5_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29539\,
            in2 => \_gnd_net_\,
            in3 => \N__27388\,
            lcout => \Lab_UT.displayAlarmZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29410\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_al_RNIHVQHE_0_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110110001"
        )
    port map (
            in0 => \N__29575\,
            in1 => \N__24084\,
            in2 => \N__24120\,
            in3 => \N__24133\,
            lcout => \Lab_UT.dictrl.nextState_al_1\,
            ltout => \Lab_UT.dictrl.nextState_al_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_al_ret_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__23571\,
            in1 => \_gnd_net_\,
            in2 => \N__23599\,
            in3 => \N__26157\,
            lcout => \Lab_UT.dictrl.un1_nextState_al24_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29410\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_al_0_0_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000111000000"
        )
    port map (
            in0 => \N__24055\,
            in1 => \N__29573\,
            in2 => \N__24127\,
            in3 => \N__23581\,
            lcout => \Lab_UT.dictrl.currState_alZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29403\,
            ce => 'H',
            sr => \N__26073\
        );

    \Lab_UT.dictrl.currState_al_0_RNIRBNK8_0_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101110111011"
        )
    port map (
            in0 => \N__24496\,
            in1 => \N__24052\,
            in2 => \N__24073\,
            in3 => \N__27355\,
            lcout => \Lab_UT.dictrl.nextState_al_1_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_0_ret_15_RNILDPC8_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000101000100"
        )
    port map (
            in0 => \N__27354\,
            in1 => \N__24068\,
            in2 => \N__23596\,
            in3 => \N__24495\,
            lcout => \Lab_UT.dictrl.nextState_al_latmux_1\,
            ltout => \Lab_UT.dictrl.nextState_al_latmux_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.nextState_al_RNISS2D9_0_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011000"
        )
    port map (
            in0 => \N__29572\,
            in1 => \N__24122\,
            in2 => \N__23575\,
            in3 => \N__24054\,
            lcout => \Lab_UT.dictrl.nextState_alZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_al_0_RNI5PG55_1_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__24056\,
            in1 => \N__27353\,
            in2 => \_gnd_net_\,
            in3 => \N__24178\,
            lcout => \Lab_UT.dictrl.N_186\,
            ltout => \Lab_UT.dictrl.N_186_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_al_0_1_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010111011"
        )
    port map (
            in0 => \N__24126\,
            in1 => \N__29574\,
            in2 => \N__24088\,
            in3 => \N__24085\,
            lcout => \Lab_UT.dictrl.currState_alZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29403\,
            ce => 'H',
            sr => \N__26073\
        );

    \Lab_UT.dictrl.currState_al_0_RNIB8DH_0_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__24072\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24053\,
            lcout => \Lab_UT.dictrl.nextState_al22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_0_ret_0_RNIHG3F_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111011101110"
        )
    port map (
            in0 => \N__23855\,
            in1 => \N__23777\,
            in2 => \N__24028\,
            in3 => \N__24013\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.un1_currState_8_u_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_ret_7_RNI03VH1_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__24886\,
            in1 => \N__24514\,
            in2 => \N__23923\,
            in3 => \N__25023\,
            lcout => \Lab_UT.dictrl.currState_ret_7_RNI03VHZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_ret_7_RNI2HHP_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24512\,
            in2 => \_gnd_net_\,
            in3 => \N__24885\,
            lcout => \Lab_UT.dictrl.un1_currState_inv_1\,
            ltout => \Lab_UT.dictrl.un1_currState_inv_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_0_ret_1_RNIPH7F1_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001100110"
        )
    port map (
            in0 => \N__23775\,
            in1 => \N__23856\,
            in2 => \N__23902\,
            in3 => \N__25021\,
            lcout => \Lab_UT.dictrl.currState_0_ret_1_RNIPH7FZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_0_ret_5_RNI9PAE_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__23869\,
            in1 => \N__23854\,
            in2 => \_gnd_net_\,
            in3 => \N__23776\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_201_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_2_RNIOB6H1_2_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23685\,
            in2 => \N__23674\,
            in3 => \N__25022\,
            lcout => \Lab_UT.dictrl.currState_2_RNIOB6H1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.r_dicRun_RNO_0_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__25024\,
            in1 => \N__24513\,
            in2 => \_gnd_net_\,
            in3 => \N__24887\,
            lcout => \Lab_UT.dictrl.r_dicRun_r_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_ret_7_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24725\,
            in2 => \_gnd_net_\,
            in3 => \N__24706\,
            lcout => \Lab_UT.dictrl.r_dicLdMtens15_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29397\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.decoder.de_atSign_4_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__24446\,
            in1 => \N__29062\,
            in2 => \N__24322\,
            in3 => \N__28539\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.decoder.de_atSignZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.decoder.de_atSign_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25225\,
            in2 => \N__24499\,
            in3 => \N__27794\,
            lcout => \Lab_UT.dictrl.de_atSign\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.decoder.de_littleA_2_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24321\,
            in3 => \N__24444\,
            lcout => \Lab_UT.dictrl.de_littleA_2\,
            ltout => \Lab_UT.dictrl.de_littleA_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.decoder.de_littleL_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__25490\,
            in1 => \N__24347\,
            in2 => \N__24484\,
            in3 => \N__27793\,
            lcout => \Lab_UT.dictrl.de_littleL\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.decoder.g0_4_2_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24445\,
            in1 => \N__24340\,
            in2 => \N__24320\,
            in3 => \N__25489\,
            lcout => \Lab_UT.dictrl.g0_4_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.decoder.de_littleN_1_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__29064\,
            in1 => \N__28756\,
            in2 => \N__24206\,
            in3 => \N__25315\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.decoder.de_littleNZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.decoder.de_littleN_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__27795\,
            in1 => \N__25402\,
            in2 => \N__25495\,
            in3 => \N__25491\,
            lcout => \Lab_UT.n_rdy\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.escKey_3_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__29063\,
            in1 => \N__28755\,
            in2 => \N__28994\,
            in3 => \N__25314\,
            lcout => \resetGen.escKeyZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_1_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28563\,
            lcout => bu_rx_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29387\,
            ce => \N__25427\,
            sr => \N__26103\
        );

    \buart.Z_rx.shifter_2_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28905\,
            lcout => bu_rx_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29387\,
            ce => \N__25427\,
            sr => \N__26103\
        );

    \Lab_UT.dictrl.decoder.de_atSign_5_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__28754\,
            in1 => \N__25376\,
            in2 => \N__28943\,
            in3 => \N__25313\,
            lcout => \Lab_UT.dictrl.decoder.de_atSignZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.uu0.l_precount_0_LC_11_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25199\,
            lcout => \Lab_UT.uu0.l_precountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29477\,
            ce => 'H',
            sr => \N__26106\
        );

    \uu2.r_addr_4_LC_11_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__25088\,
            in1 => \N__25179\,
            in2 => \_gnd_net_\,
            in3 => \N__25146\,
            lcout => \uu2.r_addrZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29473\,
            ce => 'H',
            sr => \N__26075\
        );

    \Lab_UT.displayAlarm_0_LC_11_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29548\,
            in2 => \_gnd_net_\,
            in3 => \N__27414\,
            lcout => \Lab_UT.displayAlarmZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29466\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.display.dOut_RNO_2_0_LC_11_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25867\,
            in2 => \_gnd_net_\,
            in3 => \N__25069\,
            lcout => \Lab_UT.display.N_130\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.display.dOut_RNO_0_0_LC_11_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010101110"
        )
    port map (
            in0 => \N__25659\,
            in1 => \N__25875\,
            in2 => \N__25741\,
            in3 => \N__25732\,
            lcout => OPEN,
            ltout => \Lab_UT.display.dOutP_0_iv_i_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.display.dOut_0_LC_11_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__26439\,
            in1 => \N__25708\,
            in2 => \N__25702\,
            in3 => \N__25699\,
            lcout => \L3_tx_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29466\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.displayAlarm_2_LC_11_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29547\,
            in2 => \_gnd_net_\,
            in3 => \N__27415\,
            lcout => \Lab_UT.displayAlarmZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29466\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.display.dOut_RNO_0_2_LC_11_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011001110"
        )
    port map (
            in0 => \N__25876\,
            in1 => \N__25660\,
            in2 => \N__25645\,
            in3 => \N__25633\,
            lcout => OPEN,
            ltout => \Lab_UT.display.dOutP_0_iv_i_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.display.dOut_2_LC_11_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__25816\,
            in1 => \N__26440\,
            in2 => \N__25609\,
            in3 => \N__25606\,
            lcout => \L3_tx_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29466\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.display.cnt_RNIFA8M_2_LC_11_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__26406\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26486\,
            lcout => \Lab_UT.display.un42_dOutP_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.display.cnt_RNI1STE1_1_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__25865\,
            in1 => \N__26496\,
            in2 => \_gnd_net_\,
            in3 => \N__26732\,
            lcout => \Lab_UT.display.cnt_RNI1STE1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.display.cnt_RNIE98M_2_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26401\,
            in2 => \_gnd_net_\,
            in3 => \N__26297\,
            lcout => \Lab_UT.display.N_151\,
            ltout => \Lab_UT.display.N_151_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.display.dOut_RNO_3_3_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000001010000"
        )
    port map (
            in0 => \N__26501\,
            in1 => \N__26731\,
            in2 => \N__25537\,
            in3 => \N__25534\,
            lcout => \Lab_UT.display.N_124\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.display.cnt_0_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111110"
        )
    port map (
            in0 => \N__26733\,
            in1 => \N__26402\,
            in2 => \N__26510\,
            in3 => \N__26300\,
            lcout => \Lab_UT.display.cntZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29458\,
            ce => 'H',
            sr => \N__26074\
        );

    \Lab_UT.display.cnt_2_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101011110000"
        )
    port map (
            in0 => \N__26299\,
            in1 => \_gnd_net_\,
            in2 => \N__26417\,
            in3 => \N__26500\,
            lcout => \Lab_UT.display.cntZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29458\,
            ce => 'H',
            sr => \N__26074\
        );

    \Lab_UT.display.cnt_1_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26502\,
            in2 => \_gnd_net_\,
            in3 => \N__26301\,
            lcout => \Lab_UT.display.cntZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29458\,
            ce => 'H',
            sr => \N__26074\
        );

    \Lab_UT.display.cnt_RNID88M_1_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__26298\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26495\,
            lcout => \Lab_UT.display.N_106\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.display.dOut_RNO_2_2_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25866\,
            in2 => \_gnd_net_\,
            in3 => \N__25851\,
            lcout => \Lab_UT.display.N_115\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Stens_subtractor.q_1_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__26590\,
            in1 => \N__26551\,
            in2 => \N__26960\,
            in3 => \N__26569\,
            lcout => \Lab_UT.didp.di_Stens_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29451\,
            ce => 'H',
            sr => \N__28419\
        );

    \Lab_UT.didp.Mones_subtractor.q_RNI775L5_3_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__26950\,
            in1 => \N__28024\,
            in2 => \_gnd_net_\,
            in3 => \N__27052\,
            lcout => \Lab_UT.didp.Mones_subtractor.N_80\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.display.dOut_RNO_2_1_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010100000000"
        )
    port map (
            in0 => \N__26407\,
            in1 => \N__25810\,
            in2 => \N__26334\,
            in3 => \N__26491\,
            lcout => OPEN,
            ltout => \Lab_UT.display.N_108_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.display.dOut_RNO_0_1_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011110000"
        )
    port map (
            in0 => \N__26526\,
            in1 => \N__26409\,
            in2 => \N__25783\,
            in3 => \N__25779\,
            lcout => \Lab_UT.display.dOutP_0_iv_i_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.display.cnt_RNID88M_0_1_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26490\,
            in2 => \_gnd_net_\,
            in3 => \N__26292\,
            lcout => \Lab_UT.display.N_152\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.display.cnt_RNI1STE1_2_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000001101"
        )
    port map (
            in0 => \N__26730\,
            in1 => \N__26503\,
            in2 => \N__26317\,
            in3 => \N__26410\,
            lcout => \Lab_UT.display.N_92\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.display.dOut_RNO_3_1_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__26408\,
            in1 => \N__26729\,
            in2 => \N__26365\,
            in3 => \N__26293\,
            lcout => \Lab_UT.display.N_112\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Sones_subtractor.q_RNO_0_3_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100011100001"
        )
    port map (
            in0 => \N__28197\,
            in1 => \N__26225\,
            in2 => \N__26193\,
            in3 => \N__28030\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.Sones_subtractor.q_RNO_0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Sones_subtractor.q_3_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011111010101"
        )
    port map (
            in0 => \N__28171\,
            in1 => \N__28126\,
            in2 => \N__26245\,
            in3 => \N__28996\,
            lcout => \Lab_UT.didp.di_Sones_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29443\,
            ce => 'H',
            sr => \N__28436\
        );

    \Lab_UT.didp.Sones_subtractor.q_2_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__28615\,
            in1 => \N__28125\,
            in2 => \N__26242\,
            in3 => \N__28172\,
            lcout => \Lab_UT.didp.di_Sones_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29443\,
            ce => 'H',
            sr => \N__28436\
        );

    \Lab_UT.didp.Sones_subtractor.q_RNO_0_2_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001001"
        )
    port map (
            in0 => \N__29813\,
            in1 => \N__26224\,
            in2 => \N__28102\,
            in3 => \N__28196\,
            lcout => \Lab_UT.didp.Sones_subtractor.q_RNO_0_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Sones_subtractor.q_RNIIFEO1_3_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__26223\,
            in1 => \N__28088\,
            in2 => \N__26192\,
            in3 => \N__29812\,
            lcout => \Lab_UT.didp.Sones_subtractor.un8_Mtens_ce\,
            ltout => \Lab_UT.didp.Sones_subtractor.un8_Mtens_ce_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Sones_subtractor.q_RNIP8IH2_3_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111111111"
        )
    port map (
            in0 => \N__26795\,
            in1 => \N__26760\,
            in2 => \N__26161\,
            in3 => \N__26678\,
            lcout => \Lab_UT.didp.N_82\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Sones_ce_i_0_o3_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__26679\,
            in1 => \N__26796\,
            in2 => \_gnd_net_\,
            in3 => \N__26761\,
            lcout => \Lab_UT.didp.N_81\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Sones_subtractor.q_RNIVG3M3_3_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__26713\,
            in1 => \N__26636\,
            in2 => \N__27091\,
            in3 => \N__26680\,
            lcout => \Lab_UT.didp.N_83\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Sones_subtractor.q_RNIPVIV3_3_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111111111111"
        )
    port map (
            in0 => \N__28049\,
            in1 => \N__27081\,
            in2 => \N__28021\,
            in3 => \N__26638\,
            lcout => \Lab_UT.didp.N_84\,
            ltout => \Lab_UT.didp.N_84_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Mtens_subtractor.q_RNI775L5_3_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26641\,
            in3 => \N__27046\,
            lcout => \Lab_UT.didp.q_RNI775L5_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Sones_subtractor.q_RNI0E1S4_3_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__27044\,
            in1 => \N__27085\,
            in2 => \N__28022\,
            in3 => \N__26637\,
            lcout => \Lab_UT.alarm_match\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Stens_subtractor.q_RNI775L5_3_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__28023\,
            in1 => \N__27043\,
            in2 => \N__27090\,
            in3 => \N__28161\,
            lcout => \Lab_UT.didp.Stens_subtractor.q_RNI775L5_0Z0Z_3\,
            ltout => \Lab_UT.didp.Stens_subtractor.q_RNI775L5_0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Stens_subtractor.q_RNO_1_3_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27869\,
            in2 => \N__26605\,
            in3 => \N__29701\,
            lcout => \Lab_UT.didp.Stens_subtractor.un1_q_c2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Sones_subtractor.q_RNI775L5_3_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28050\,
            in2 => \_gnd_net_\,
            in3 => \N__27345\,
            lcout => \Lab_UT.didp.Sones_subtractor.q_RNI775L5_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Stens_subtractor.q_RNO_0_1_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010111000101"
        )
    port map (
            in0 => \N__26583\,
            in1 => \N__26565\,
            in2 => \N__28175\,
            in3 => \N__28818\,
            lcout => \Lab_UT.didp.Stens_subtractor.q_7_i_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Mtens_subtractor.q_RNO_2_1_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100001"
        )
    port map (
            in0 => \N__28684\,
            in1 => \N__30030\,
            in2 => \N__27949\,
            in3 => \N__27045\,
            lcout => \Lab_UT.didp.Mtens_subtractor.q_RNO_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Mtens_subtractor.q_RNO_0_2_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010011100"
        )
    port map (
            in0 => \N__30028\,
            in1 => \N__26872\,
            in2 => \N__26899\,
            in3 => \N__27943\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.Mtens_subtractor.q_RNO_0_3_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Mtens_subtractor.q_2_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110111101100"
        )
    port map (
            in0 => \N__27981\,
            in1 => \N__26919\,
            in2 => \N__26974\,
            in3 => \N__28614\,
            lcout => \Lab_UT.di_Mtens_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29429\,
            ce => 'H',
            sr => \N__28446\
        );

    \Lab_UT.didp.Mtens_subtractor.q_RNIE7IL1_3_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__30027\,
            in1 => \N__26870\,
            in2 => \N__26831\,
            in3 => \N__27942\,
            lcout => \Lab_UT.didp.un3_Mtens_rst\,
            ltout => \Lab_UT.didp.un3_Mtens_rst_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Mtens_subtractor.q_RNO_0_0_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110100000010"
        )
    port map (
            in0 => \N__28020\,
            in1 => \N__26961\,
            in2 => \N__26932\,
            in3 => \N__30029\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.Mtens_subtractor.un1_q_axb0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Mtens_subtractor.q_0_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101111101010"
        )
    port map (
            in0 => \N__26918\,
            in1 => \N__27980\,
            in2 => \N__26902\,
            in3 => \N__29097\,
            lcout => \Lab_UT.didp.di_MtensZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29429\,
            ce => 'H',
            sr => \N__28446\
        );

    \Lab_UT.didp.Stens_subtractor.q_RNI775L5_0_3_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__28019\,
            in1 => \N__27050\,
            in2 => \N__27089\,
            in3 => \N__28179\,
            lcout => \Lab_UT.didp.Mtens_ce\,
            ltout => \Lab_UT.didp.Mtens_ce_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Mtens_subtractor.q_RNO_0_3_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010011010011010"
        )
    port map (
            in0 => \N__26824\,
            in1 => \N__26871\,
            in2 => \N__26839\,
            in3 => \N__27958\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.Mtens_subtractor.q_RNO_0_2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Mtens_subtractor.q_3_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__27982\,
            in1 => \_gnd_net_\,
            in2 => \N__26836\,
            in3 => \N__28987\,
            lcout => \Lab_UT.didp.di_Mtens_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29429\,
            ce => 'H',
            sr => \N__28446\
        );

    \Lab_UT.didp.Mones_subtractor.q_RNIN8C59_3_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010010000000"
        )
    port map (
            in0 => \N__29950\,
            in1 => \N__30107\,
            in2 => \N__27325\,
            in3 => \N__27435\,
            lcout => \Lab_UT.didp.Mones_subtractor.q_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.dicLdMones_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101011001100"
        )
    port map (
            in0 => \N__27436\,
            in1 => \N__27324\,
            in2 => \N__29962\,
            in3 => \N__29891\,
            lcout => \Lab_UT.dicLdMones\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29420\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.dicLdMtens_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__29892\,
            in1 => \N__27006\,
            in2 => \N__26992\,
            in3 => \N__29956\,
            lcout => \Lab_UT.dicLdMtens\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29420\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_0_ret_6_RNIU5JA3_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__27313\,
            in1 => \N__27813\,
            in2 => \_gnd_net_\,
            in3 => \N__27301\,
            lcout => \Lab_UT.dicLdMtens_latmux\,
            ltout => \Lab_UT.dicLdMtens_latmux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Mtens_subtractor.q_7_i_o2_2_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011111111111"
        )
    port map (
            in0 => \N__29951\,
            in1 => \N__27002\,
            in2 => \N__27169\,
            in3 => \N__28682\,
            lcout => \Lab_UT.didp.Mtens_subtractor.N_87\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Stens_subtractor.q_RNI68H41_3_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__27166\,
            in1 => \N__27870\,
            in2 => \N__27130\,
            in3 => \N__29699\,
            lcout => \Lab_UT.didp.un6_Mtens_ce\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Mtens_subtractor.q_RNO_0_1_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010111110"
        )
    port map (
            in0 => \N__27051\,
            in1 => \N__30037\,
            in2 => \N__27947\,
            in3 => \N__28683\,
            lcout => \Lab_UT.didp.Mtens_subtractor.N_145\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Mtens_subtractor.q_RNO_1_1_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000010011"
        )
    port map (
            in0 => \N__29952\,
            in1 => \N__27016\,
            in2 => \N__27007\,
            in3 => \N__26988\,
            lcout => \Lab_UT.didp.Mtens_subtractor.N_147\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Mtens_subtractor.q_1_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001010100"
        )
    port map (
            in0 => \N__26980\,
            in1 => \N__27979\,
            in2 => \N__28822\,
            in3 => \N__27964\,
            lcout => \Lab_UT.didp.di_Mtens_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29412\,
            ce => 'H',
            sr => \N__28456\
        );

    \Lab_UT.didp.Mtens_subtractor.q_RNO_1_3_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__28678\,
            in1 => \N__30039\,
            in2 => \_gnd_net_\,
            in3 => \N__27934\,
            lcout => \Lab_UT.didp.Mtens_subtractor.un1_q_c2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Mones_subtractor.q_RNITOVP_1_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__30081\,
            in1 => \N__27938\,
            in2 => \_gnd_net_\,
            in3 => \N__29780\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.q_RNITOVP_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.curr_LED_RNIJFM52_1_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__27832\,
            in1 => \_gnd_net_\,
            in2 => \N__27892\,
            in3 => \N__29644\,
            lcout => led_c_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Stens_subtractor.q_RNI99F11_1_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__27871\,
            in1 => \N__29781\,
            in2 => \_gnd_net_\,
            in3 => \N__28105\,
            lcout => \Lab_UT.didp.q_RNI99F11_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.currState_0_ret_12_RNIB2D93_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__27826\,
            in1 => \N__27812\,
            in2 => \_gnd_net_\,
            in3 => \N__27562\,
            lcout => \Lab_UT.dicLdMones_latmux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.displayAlarm_6_LC_12_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29532\,
            lcout => \Lab_UT.displayAlarmZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29474\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.displayAlarm_4_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29546\,
            in2 => \_gnd_net_\,
            in3 => \N__27413\,
            lcout => \Lab_UT.displayAlarmZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29467\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Sones_subtractor.q_RNO_1_1_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001001"
        )
    port map (
            in0 => \N__27341\,
            in1 => \N__28092\,
            in2 => \N__28059\,
            in3 => \N__29814\,
            lcout => \Lab_UT.didp.Sones_subtractor.q_RNO_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.dicLdSones_RNISPBP3_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__29961\,
            in1 => \_gnd_net_\,
            in2 => \N__29845\,
            in3 => \N__29867\,
            lcout => OPEN,
            ltout => \Lab_UT.ld_enable_Sones_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Sones_subtractor.q_RNO_0_1_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001011111"
        )
    port map (
            in0 => \N__28055\,
            in1 => \_gnd_net_\,
            in2 => \N__28210\,
            in3 => \N__28207\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.Sones_subtractor.q_7_i_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Sones_subtractor.q_1_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000001000"
        )
    port map (
            in0 => \N__28124\,
            in1 => \N__28174\,
            in2 => \N__28201\,
            in3 => \N__28820\,
            lcout => \Lab_UT.didp.di_Sones_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29452\,
            ce => 'H',
            sr => \N__28455\
        );

    \Lab_UT.didp.Sones_subtractor.q_RNO_0_0_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28198\,
            in2 => \_gnd_net_\,
            in3 => \N__29816\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.Sones_subtractor.un1_q_axb0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Sones_subtractor.q_0_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110110011"
        )
    port map (
            in0 => \N__28123\,
            in1 => \N__28173\,
            in2 => \N__28129\,
            in3 => \N__29107\,
            lcout => \Lab_UT.didp.di_Sones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29452\,
            ce => 'H',
            sr => \N__28455\
        );

    \Lab_UT.didp.Sones_subtractor.q_7_i_o2_3_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111101011111"
        )
    port map (
            in0 => \N__29868\,
            in1 => \N__29843\,
            in2 => \N__28060\,
            in3 => \N__29960\,
            lcout => \Lab_UT.didp.Sones_subtractor.N_85\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Sones_subtractor.q_RNO_1_3_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111010"
        )
    port map (
            in0 => \N__29815\,
            in1 => \_gnd_net_\,
            in2 => \N__28103\,
            in3 => \N__28051\,
            lcout => \Lab_UT.didp.Sones_subtractor.un1_q_c2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Mones_subtractor.q_RNIQEF9_3_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__28285\,
            in1 => \N__30072\,
            in2 => \N__28247\,
            in3 => \N__29985\,
            lcout => \Lab_UT.didp.un4_Mtens_ce\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Mones_subtractor.q_RNO_0_0_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__29986\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30120\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.Mones_subtractor.un1_q_axb_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Mones_subtractor.q_0_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110101110101"
        )
    port map (
            in0 => \N__28660\,
            in1 => \N__28633\,
            in2 => \N__29110\,
            in3 => \N__29098\,
            lcout => \Lab_UT.didp.di_Mones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29444\,
            ce => 'H',
            sr => \N__28447\
        );

    \Lab_UT.didp.Mones_subtractor.q_3_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101110011"
        )
    port map (
            in0 => \N__28636\,
            in1 => \N__28665\,
            in2 => \N__30136\,
            in3 => \N__28980\,
            lcout => \Lab_UT.didp.di_Mones_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29444\,
            ce => 'H',
            sr => \N__28447\
        );

    \Lab_UT.didp.Mones_subtractor.q_1_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110000000100000"
        )
    port map (
            in0 => \N__30046\,
            in1 => \N__28634\,
            in2 => \N__28677\,
            in3 => \N__28819\,
            lcout => \Lab_UT.didp.di_Mones_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29444\,
            ce => 'H',
            sr => \N__28447\
        );

    \Lab_UT.didp.Mones_subtractor.q_RNO_0_2_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000010001"
        )
    port map (
            in0 => \N__28264\,
            in1 => \N__30121\,
            in2 => \_gnd_net_\,
            in3 => \N__28286\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.Mones_subtractor.q_RNO_0_2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Mones_subtractor.q_2_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100000100000"
        )
    port map (
            in0 => \N__28664\,
            in1 => \N__28635\,
            in2 => \N__28618\,
            in3 => \N__28607\,
            lcout => \Lab_UT.didp.di_Mones_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29444\,
            ce => 'H',
            sr => \N__28447\
        );

    \Lab_UT.didp.Mones_subtractor.un1_q_cry_0_s1_c_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29987\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_9_0_\,
            carryout => \Lab_UT.didp.Mones_subtractor.un1_q_cry_0_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Mones_subtractor.un1_q_cry_0_s1_THRU_LUT4_0_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30073\,
            in2 => \N__28357\,
            in3 => \N__28360\,
            lcout => \Lab_UT.didp.Mones_subtractor.un1_q_cry_0_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \Lab_UT.didp.Mones_subtractor.un1_q_cry_0_s1\,
            carryout => \Lab_UT.didp.Mones_subtractor.un1_q_cry_1_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Mones_subtractor.un1_q_cry_1_s1_THRU_LUT4_0_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28353\,
            in2 => \N__28295\,
            in3 => \N__28255\,
            lcout => \Lab_UT.didp.Mones_subtractor.un1_q_cry_1_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \Lab_UT.didp.Mones_subtractor.un1_q_cry_1_s1\,
            carryout => \Lab_UT.didp.Mones_subtractor.un1_q_cry_2_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Mones_subtractor.q_RNO_0_3_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010011001"
        )
    port map (
            in0 => \N__28240\,
            in1 => \N__30119\,
            in2 => \_gnd_net_\,
            in3 => \N__28213\,
            lcout => \Lab_UT.didp.Mones_subtractor.q_RNO_0_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Mones_subtractor.q_RNO_0_1_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000010001"
        )
    port map (
            in0 => \N__30127\,
            in1 => \N__30118\,
            in2 => \_gnd_net_\,
            in3 => \N__30074\,
            lcout => \Lab_UT.didp.Mones_subtractor.q_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Mones_subtractor.q_RNIRMVP_0_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__30040\,
            in1 => \N__29774\,
            in2 => \_gnd_net_\,
            in3 => \N__29988\,
            lcout => \Lab_UT.didp.q_RNIRMVP_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.dicLdSones_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__29957\,
            in1 => \N__29893\,
            in2 => \N__29844\,
            in3 => \N__29869\,
            lcout => \Lab_UT.dicLdSones\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29430\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.Stens_subtractor.q_RNI77F11_0_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__29821\,
            in1 => \N__29782\,
            in2 => \_gnd_net_\,
            in3 => \N__29700\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.q_RNI77F11_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.curr_LED_RNIFBM52_1_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29653\,
            in2 => \N__29647\,
            in3 => \N__29637\,
            lcout => led_c_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.r_dicAlarmIdle_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29512\,
            in2 => \_gnd_net_\,
            in3 => \N__29584\,
            lcout => \Lab_UT.alarm_off\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29421\,
            ce => 'H',
            sr => \N__29131\
        );
end \INTERFACE\;
