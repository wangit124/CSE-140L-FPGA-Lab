// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     Jun 5 2019 04:46:17

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "latticehx1k" view "INTERFACE"

module latticehx1k (
    led,
    o_serial_data,
    to_ir,
    sd,
    from_pc,
    clk_in);

    output [4:0] led;
    output o_serial_data;
    output to_ir;
    output sd;
    input from_pc;
    input clk_in;

    wire N__30236;
    wire N__30235;
    wire N__30234;
    wire N__30227;
    wire N__30226;
    wire N__30225;
    wire N__30218;
    wire N__30217;
    wire N__30216;
    wire N__30209;
    wire N__30208;
    wire N__30207;
    wire N__30200;
    wire N__30199;
    wire N__30198;
    wire N__30191;
    wire N__30190;
    wire N__30189;
    wire N__30182;
    wire N__30181;
    wire N__30180;
    wire N__30173;
    wire N__30172;
    wire N__30171;
    wire N__30164;
    wire N__30163;
    wire N__30162;
    wire N__30155;
    wire N__30154;
    wire N__30153;
    wire N__30136;
    wire N__30133;
    wire N__30130;
    wire N__30127;
    wire N__30124;
    wire N__30121;
    wire N__30120;
    wire N__30119;
    wire N__30118;
    wire N__30113;
    wire N__30108;
    wire N__30107;
    wire N__30104;
    wire N__30101;
    wire N__30098;
    wire N__30095;
    wire N__30092;
    wire N__30089;
    wire N__30082;
    wire N__30081;
    wire N__30078;
    wire N__30075;
    wire N__30074;
    wire N__30073;
    wire N__30072;
    wire N__30069;
    wire N__30066;
    wire N__30061;
    wire N__30058;
    wire N__30055;
    wire N__30046;
    wire N__30043;
    wire N__30040;
    wire N__30039;
    wire N__30038;
    wire N__30037;
    wire N__30034;
    wire N__30031;
    wire N__30030;
    wire N__30029;
    wire N__30028;
    wire N__30027;
    wire N__30024;
    wire N__30021;
    wire N__30016;
    wire N__30013;
    wire N__30006;
    wire N__30003;
    wire N__29992;
    wire N__29989;
    wire N__29988;
    wire N__29987;
    wire N__29986;
    wire N__29985;
    wire N__29982;
    wire N__29977;
    wire N__29972;
    wire N__29969;
    wire N__29962;
    wire N__29961;
    wire N__29960;
    wire N__29959;
    wire N__29958;
    wire N__29957;
    wire N__29956;
    wire N__29953;
    wire N__29952;
    wire N__29951;
    wire N__29950;
    wire N__29945;
    wire N__29940;
    wire N__29939;
    wire N__29936;
    wire N__29929;
    wire N__29924;
    wire N__29921;
    wire N__29918;
    wire N__29915;
    wire N__29912;
    wire N__29905;
    wire N__29902;
    wire N__29893;
    wire N__29892;
    wire N__29891;
    wire N__29888;
    wire N__29883;
    wire N__29882;
    wire N__29877;
    wire N__29874;
    wire N__29869;
    wire N__29868;
    wire N__29867;
    wire N__29864;
    wire N__29859;
    wire N__29854;
    wire N__29851;
    wire N__29848;
    wire N__29845;
    wire N__29844;
    wire N__29843;
    wire N__29840;
    wire N__29837;
    wire N__29832;
    wire N__29829;
    wire N__29826;
    wire N__29821;
    wire N__29820;
    wire N__29817;
    wire N__29816;
    wire N__29815;
    wire N__29814;
    wire N__29813;
    wire N__29812;
    wire N__29809;
    wire N__29806;
    wire N__29799;
    wire N__29794;
    wire N__29791;
    wire N__29782;
    wire N__29781;
    wire N__29780;
    wire N__29779;
    wire N__29778;
    wire N__29775;
    wire N__29774;
    wire N__29773;
    wire N__29768;
    wire N__29765;
    wire N__29762;
    wire N__29761;
    wire N__29758;
    wire N__29755;
    wire N__29752;
    wire N__29749;
    wire N__29744;
    wire N__29741;
    wire N__29736;
    wire N__29733;
    wire N__29726;
    wire N__29725;
    wire N__29724;
    wire N__29721;
    wire N__29718;
    wire N__29715;
    wire N__29710;
    wire N__29701;
    wire N__29700;
    wire N__29699;
    wire N__29696;
    wire N__29693;
    wire N__29690;
    wire N__29689;
    wire N__29686;
    wire N__29685;
    wire N__29684;
    wire N__29683;
    wire N__29678;
    wire N__29675;
    wire N__29672;
    wire N__29665;
    wire N__29660;
    wire N__29653;
    wire N__29650;
    wire N__29647;
    wire N__29644;
    wire N__29641;
    wire N__29638;
    wire N__29637;
    wire N__29634;
    wire N__29631;
    wire N__29630;
    wire N__29629;
    wire N__29624;
    wire N__29619;
    wire N__29616;
    wire N__29613;
    wire N__29612;
    wire N__29609;
    wire N__29606;
    wire N__29603;
    wire N__29596;
    wire N__29593;
    wire N__29590;
    wire N__29587;
    wire N__29584;
    wire N__29581;
    wire N__29578;
    wire N__29577;
    wire N__29576;
    wire N__29575;
    wire N__29574;
    wire N__29573;
    wire N__29572;
    wire N__29569;
    wire N__29562;
    wire N__29555;
    wire N__29548;
    wire N__29547;
    wire N__29546;
    wire N__29541;
    wire N__29540;
    wire N__29539;
    wire N__29536;
    wire N__29533;
    wire N__29532;
    wire N__29529;
    wire N__29526;
    wire N__29521;
    wire N__29518;
    wire N__29513;
    wire N__29512;
    wire N__29509;
    wire N__29506;
    wire N__29503;
    wire N__29500;
    wire N__29491;
    wire N__29490;
    wire N__29487;
    wire N__29484;
    wire N__29481;
    wire N__29480;
    wire N__29479;
    wire N__29478;
    wire N__29477;
    wire N__29476;
    wire N__29475;
    wire N__29474;
    wire N__29473;
    wire N__29472;
    wire N__29471;
    wire N__29470;
    wire N__29469;
    wire N__29468;
    wire N__29467;
    wire N__29466;
    wire N__29465;
    wire N__29464;
    wire N__29463;
    wire N__29462;
    wire N__29461;
    wire N__29460;
    wire N__29459;
    wire N__29458;
    wire N__29457;
    wire N__29456;
    wire N__29455;
    wire N__29454;
    wire N__29453;
    wire N__29452;
    wire N__29451;
    wire N__29450;
    wire N__29449;
    wire N__29448;
    wire N__29447;
    wire N__29446;
    wire N__29445;
    wire N__29444;
    wire N__29443;
    wire N__29442;
    wire N__29441;
    wire N__29440;
    wire N__29439;
    wire N__29438;
    wire N__29437;
    wire N__29436;
    wire N__29435;
    wire N__29434;
    wire N__29433;
    wire N__29432;
    wire N__29431;
    wire N__29430;
    wire N__29429;
    wire N__29428;
    wire N__29427;
    wire N__29426;
    wire N__29425;
    wire N__29424;
    wire N__29423;
    wire N__29422;
    wire N__29421;
    wire N__29420;
    wire N__29419;
    wire N__29418;
    wire N__29417;
    wire N__29416;
    wire N__29415;
    wire N__29414;
    wire N__29413;
    wire N__29412;
    wire N__29411;
    wire N__29410;
    wire N__29409;
    wire N__29408;
    wire N__29407;
    wire N__29406;
    wire N__29405;
    wire N__29404;
    wire N__29403;
    wire N__29402;
    wire N__29401;
    wire N__29400;
    wire N__29399;
    wire N__29398;
    wire N__29397;
    wire N__29396;
    wire N__29395;
    wire N__29394;
    wire N__29393;
    wire N__29392;
    wire N__29391;
    wire N__29390;
    wire N__29389;
    wire N__29388;
    wire N__29387;
    wire N__29386;
    wire N__29385;
    wire N__29384;
    wire N__29383;
    wire N__29382;
    wire N__29381;
    wire N__29380;
    wire N__29379;
    wire N__29378;
    wire N__29377;
    wire N__29376;
    wire N__29375;
    wire N__29374;
    wire N__29373;
    wire N__29372;
    wire N__29371;
    wire N__29370;
    wire N__29367;
    wire N__29364;
    wire N__29137;
    wire N__29134;
    wire N__29131;
    wire N__29130;
    wire N__29127;
    wire N__29126;
    wire N__29123;
    wire N__29120;
    wire N__29115;
    wire N__29110;
    wire N__29107;
    wire N__29106;
    wire N__29105;
    wire N__29104;
    wire N__29103;
    wire N__29102;
    wire N__29099;
    wire N__29098;
    wire N__29097;
    wire N__29094;
    wire N__29091;
    wire N__29086;
    wire N__29083;
    wire N__29080;
    wire N__29077;
    wire N__29074;
    wire N__29073;
    wire N__29070;
    wire N__29065;
    wire N__29064;
    wire N__29063;
    wire N__29062;
    wire N__29059;
    wire N__29052;
    wire N__29049;
    wire N__29048;
    wire N__29047;
    wire N__29042;
    wire N__29035;
    wire N__29030;
    wire N__29027;
    wire N__29026;
    wire N__29023;
    wire N__29020;
    wire N__29015;
    wire N__29010;
    wire N__29003;
    wire N__28996;
    wire N__28995;
    wire N__28994;
    wire N__28991;
    wire N__28988;
    wire N__28987;
    wire N__28986;
    wire N__28985;
    wire N__28984;
    wire N__28983;
    wire N__28982;
    wire N__28981;
    wire N__28980;
    wire N__28979;
    wire N__28978;
    wire N__28975;
    wire N__28974;
    wire N__28971;
    wire N__28968;
    wire N__28965;
    wire N__28964;
    wire N__28957;
    wire N__28954;
    wire N__28951;
    wire N__28948;
    wire N__28947;
    wire N__28944;
    wire N__28943;
    wire N__28938;
    wire N__28935;
    wire N__28932;
    wire N__28925;
    wire N__28924;
    wire N__28921;
    wire N__28916;
    wire N__28913;
    wire N__28910;
    wire N__28907;
    wire N__28906;
    wire N__28905;
    wire N__28902;
    wire N__28899;
    wire N__28896;
    wire N__28893;
    wire N__28890;
    wire N__28887;
    wire N__28884;
    wire N__28881;
    wire N__28878;
    wire N__28873;
    wire N__28870;
    wire N__28867;
    wire N__28864;
    wire N__28861;
    wire N__28858;
    wire N__28851;
    wire N__28844;
    wire N__28837;
    wire N__28822;
    wire N__28821;
    wire N__28820;
    wire N__28819;
    wire N__28818;
    wire N__28817;
    wire N__28816;
    wire N__28813;
    wire N__28812;
    wire N__28809;
    wire N__28806;
    wire N__28803;
    wire N__28800;
    wire N__28797;
    wire N__28796;
    wire N__28795;
    wire N__28792;
    wire N__28789;
    wire N__28786;
    wire N__28783;
    wire N__28776;
    wire N__28773;
    wire N__28772;
    wire N__28771;
    wire N__28766;
    wire N__28763;
    wire N__28760;
    wire N__28757;
    wire N__28756;
    wire N__28755;
    wire N__28754;
    wire N__28753;
    wire N__28750;
    wire N__28747;
    wire N__28744;
    wire N__28743;
    wire N__28738;
    wire N__28735;
    wire N__28732;
    wire N__28729;
    wire N__28726;
    wire N__28721;
    wire N__28718;
    wire N__28715;
    wire N__28708;
    wire N__28705;
    wire N__28684;
    wire N__28683;
    wire N__28682;
    wire N__28679;
    wire N__28678;
    wire N__28677;
    wire N__28672;
    wire N__28669;
    wire N__28666;
    wire N__28665;
    wire N__28664;
    wire N__28661;
    wire N__28660;
    wire N__28653;
    wire N__28644;
    wire N__28641;
    wire N__28636;
    wire N__28635;
    wire N__28634;
    wire N__28633;
    wire N__28624;
    wire N__28621;
    wire N__28618;
    wire N__28615;
    wire N__28614;
    wire N__28613;
    wire N__28612;
    wire N__28611;
    wire N__28610;
    wire N__28609;
    wire N__28608;
    wire N__28607;
    wire N__28606;
    wire N__28603;
    wire N__28602;
    wire N__28601;
    wire N__28598;
    wire N__28597;
    wire N__28596;
    wire N__28593;
    wire N__28590;
    wire N__28585;
    wire N__28580;
    wire N__28577;
    wire N__28574;
    wire N__28573;
    wire N__28570;
    wire N__28567;
    wire N__28564;
    wire N__28563;
    wire N__28560;
    wire N__28557;
    wire N__28554;
    wire N__28551;
    wire N__28548;
    wire N__28543;
    wire N__28540;
    wire N__28539;
    wire N__28536;
    wire N__28533;
    wire N__28530;
    wire N__28527;
    wire N__28524;
    wire N__28521;
    wire N__28518;
    wire N__28515;
    wire N__28510;
    wire N__28509;
    wire N__28508;
    wire N__28507;
    wire N__28500;
    wire N__28497;
    wire N__28494;
    wire N__28485;
    wire N__28476;
    wire N__28469;
    wire N__28456;
    wire N__28455;
    wire N__28452;
    wire N__28449;
    wire N__28448;
    wire N__28447;
    wire N__28446;
    wire N__28443;
    wire N__28440;
    wire N__28437;
    wire N__28436;
    wire N__28433;
    wire N__28430;
    wire N__28423;
    wire N__28420;
    wire N__28419;
    wire N__28416;
    wire N__28413;
    wire N__28408;
    wire N__28405;
    wire N__28402;
    wire N__28399;
    wire N__28396;
    wire N__28393;
    wire N__28390;
    wire N__28387;
    wire N__28384;
    wire N__28381;
    wire N__28378;
    wire N__28375;
    wire N__28372;
    wire N__28369;
    wire N__28360;
    wire N__28357;
    wire N__28356;
    wire N__28355;
    wire N__28354;
    wire N__28353;
    wire N__28350;
    wire N__28347;
    wire N__28344;
    wire N__28341;
    wire N__28336;
    wire N__28333;
    wire N__28330;
    wire N__28327;
    wire N__28324;
    wire N__28321;
    wire N__28318;
    wire N__28315;
    wire N__28312;
    wire N__28309;
    wire N__28304;
    wire N__28297;
    wire N__28296;
    wire N__28295;
    wire N__28290;
    wire N__28287;
    wire N__28286;
    wire N__28285;
    wire N__28282;
    wire N__28279;
    wire N__28274;
    wire N__28271;
    wire N__28264;
    wire N__28261;
    wire N__28258;
    wire N__28255;
    wire N__28252;
    wire N__28251;
    wire N__28248;
    wire N__28247;
    wire N__28244;
    wire N__28241;
    wire N__28240;
    wire N__28237;
    wire N__28234;
    wire N__28231;
    wire N__28228;
    wire N__28225;
    wire N__28222;
    wire N__28213;
    wire N__28210;
    wire N__28207;
    wire N__28204;
    wire N__28201;
    wire N__28198;
    wire N__28197;
    wire N__28196;
    wire N__28193;
    wire N__28188;
    wire N__28185;
    wire N__28180;
    wire N__28179;
    wire N__28176;
    wire N__28175;
    wire N__28174;
    wire N__28173;
    wire N__28172;
    wire N__28171;
    wire N__28168;
    wire N__28165;
    wire N__28162;
    wire N__28161;
    wire N__28156;
    wire N__28151;
    wire N__28148;
    wire N__28145;
    wire N__28140;
    wire N__28129;
    wire N__28126;
    wire N__28125;
    wire N__28124;
    wire N__28123;
    wire N__28120;
    wire N__28117;
    wire N__28112;
    wire N__28105;
    wire N__28104;
    wire N__28103;
    wire N__28102;
    wire N__28099;
    wire N__28096;
    wire N__28093;
    wire N__28092;
    wire N__28089;
    wire N__28088;
    wire N__28085;
    wire N__28082;
    wire N__28077;
    wire N__28072;
    wire N__28067;
    wire N__28060;
    wire N__28059;
    wire N__28056;
    wire N__28055;
    wire N__28052;
    wire N__28051;
    wire N__28050;
    wire N__28049;
    wire N__28040;
    wire N__28035;
    wire N__28030;
    wire N__28027;
    wire N__28024;
    wire N__28023;
    wire N__28022;
    wire N__28021;
    wire N__28020;
    wire N__28019;
    wire N__28016;
    wire N__28013;
    wire N__28010;
    wire N__28007;
    wire N__28002;
    wire N__27999;
    wire N__27996;
    wire N__27991;
    wire N__27982;
    wire N__27981;
    wire N__27980;
    wire N__27979;
    wire N__27972;
    wire N__27969;
    wire N__27964;
    wire N__27961;
    wire N__27958;
    wire N__27955;
    wire N__27952;
    wire N__27949;
    wire N__27948;
    wire N__27947;
    wire N__27944;
    wire N__27943;
    wire N__27942;
    wire N__27939;
    wire N__27938;
    wire N__27935;
    wire N__27934;
    wire N__27931;
    wire N__27926;
    wire N__27923;
    wire N__27920;
    wire N__27917;
    wire N__27914;
    wire N__27911;
    wire N__27908;
    wire N__27905;
    wire N__27892;
    wire N__27889;
    wire N__27886;
    wire N__27883;
    wire N__27880;
    wire N__27877;
    wire N__27874;
    wire N__27873;
    wire N__27872;
    wire N__27871;
    wire N__27870;
    wire N__27869;
    wire N__27864;
    wire N__27861;
    wire N__27858;
    wire N__27855;
    wire N__27852;
    wire N__27847;
    wire N__27842;
    wire N__27837;
    wire N__27832;
    wire N__27829;
    wire N__27826;
    wire N__27823;
    wire N__27820;
    wire N__27817;
    wire N__27814;
    wire N__27813;
    wire N__27812;
    wire N__27811;
    wire N__27810;
    wire N__27809;
    wire N__27808;
    wire N__27807;
    wire N__27806;
    wire N__27803;
    wire N__27802;
    wire N__27799;
    wire N__27796;
    wire N__27795;
    wire N__27794;
    wire N__27793;
    wire N__27792;
    wire N__27791;
    wire N__27790;
    wire N__27789;
    wire N__27788;
    wire N__27787;
    wire N__27784;
    wire N__27783;
    wire N__27782;
    wire N__27781;
    wire N__27778;
    wire N__27777;
    wire N__27774;
    wire N__27773;
    wire N__27766;
    wire N__27761;
    wire N__27756;
    wire N__27749;
    wire N__27748;
    wire N__27747;
    wire N__27746;
    wire N__27745;
    wire N__27740;
    wire N__27735;
    wire N__27732;
    wire N__27731;
    wire N__27730;
    wire N__27729;
    wire N__27726;
    wire N__27725;
    wire N__27722;
    wire N__27717;
    wire N__27716;
    wire N__27713;
    wire N__27712;
    wire N__27711;
    wire N__27710;
    wire N__27705;
    wire N__27702;
    wire N__27701;
    wire N__27700;
    wire N__27697;
    wire N__27692;
    wire N__27687;
    wire N__27684;
    wire N__27677;
    wire N__27672;
    wire N__27665;
    wire N__27662;
    wire N__27659;
    wire N__27656;
    wire N__27651;
    wire N__27648;
    wire N__27647;
    wire N__27646;
    wire N__27645;
    wire N__27644;
    wire N__27643;
    wire N__27640;
    wire N__27637;
    wire N__27632;
    wire N__27629;
    wire N__27626;
    wire N__27621;
    wire N__27612;
    wire N__27605;
    wire N__27594;
    wire N__27583;
    wire N__27562;
    wire N__27561;
    wire N__27560;
    wire N__27559;
    wire N__27556;
    wire N__27553;
    wire N__27552;
    wire N__27551;
    wire N__27546;
    wire N__27545;
    wire N__27544;
    wire N__27543;
    wire N__27542;
    wire N__27541;
    wire N__27538;
    wire N__27535;
    wire N__27532;
    wire N__27529;
    wire N__27526;
    wire N__27521;
    wire N__27518;
    wire N__27517;
    wire N__27512;
    wire N__27511;
    wire N__27510;
    wire N__27507;
    wire N__27504;
    wire N__27501;
    wire N__27498;
    wire N__27493;
    wire N__27490;
    wire N__27487;
    wire N__27484;
    wire N__27483;
    wire N__27482;
    wire N__27479;
    wire N__27476;
    wire N__27475;
    wire N__27468;
    wire N__27461;
    wire N__27456;
    wire N__27445;
    wire N__27436;
    wire N__27435;
    wire N__27430;
    wire N__27427;
    wire N__27424;
    wire N__27421;
    wire N__27418;
    wire N__27415;
    wire N__27414;
    wire N__27413;
    wire N__27408;
    wire N__27405;
    wire N__27402;
    wire N__27399;
    wire N__27396;
    wire N__27395;
    wire N__27392;
    wire N__27389;
    wire N__27388;
    wire N__27385;
    wire N__27382;
    wire N__27379;
    wire N__27374;
    wire N__27367;
    wire N__27364;
    wire N__27361;
    wire N__27358;
    wire N__27355;
    wire N__27354;
    wire N__27353;
    wire N__27346;
    wire N__27345;
    wire N__27342;
    wire N__27341;
    wire N__27338;
    wire N__27335;
    wire N__27332;
    wire N__27325;
    wire N__27324;
    wire N__27321;
    wire N__27316;
    wire N__27313;
    wire N__27310;
    wire N__27307;
    wire N__27304;
    wire N__27301;
    wire N__27300;
    wire N__27299;
    wire N__27298;
    wire N__27297;
    wire N__27296;
    wire N__27295;
    wire N__27294;
    wire N__27293;
    wire N__27292;
    wire N__27289;
    wire N__27286;
    wire N__27285;
    wire N__27284;
    wire N__27281;
    wire N__27278;
    wire N__27277;
    wire N__27276;
    wire N__27271;
    wire N__27264;
    wire N__27261;
    wire N__27258;
    wire N__27255;
    wire N__27250;
    wire N__27249;
    wire N__27248;
    wire N__27247;
    wire N__27246;
    wire N__27243;
    wire N__27240;
    wire N__27235;
    wire N__27232;
    wire N__27227;
    wire N__27220;
    wire N__27213;
    wire N__27212;
    wire N__27211;
    wire N__27210;
    wire N__27209;
    wire N__27206;
    wire N__27201;
    wire N__27194;
    wire N__27189;
    wire N__27180;
    wire N__27169;
    wire N__27166;
    wire N__27163;
    wire N__27162;
    wire N__27161;
    wire N__27160;
    wire N__27159;
    wire N__27156;
    wire N__27153;
    wire N__27148;
    wire N__27145;
    wire N__27142;
    wire N__27139;
    wire N__27130;
    wire N__27127;
    wire N__27126;
    wire N__27123;
    wire N__27120;
    wire N__27119;
    wire N__27118;
    wire N__27115;
    wire N__27112;
    wire N__27109;
    wire N__27106;
    wire N__27103;
    wire N__27100;
    wire N__27091;
    wire N__27090;
    wire N__27089;
    wire N__27086;
    wire N__27085;
    wire N__27082;
    wire N__27081;
    wire N__27078;
    wire N__27075;
    wire N__27068;
    wire N__27065;
    wire N__27062;
    wire N__27059;
    wire N__27052;
    wire N__27051;
    wire N__27050;
    wire N__27047;
    wire N__27046;
    wire N__27045;
    wire N__27044;
    wire N__27043;
    wire N__27040;
    wire N__27037;
    wire N__27034;
    wire N__27025;
    wire N__27016;
    wire N__27013;
    wire N__27010;
    wire N__27007;
    wire N__27006;
    wire N__27003;
    wire N__27002;
    wire N__26995;
    wire N__26992;
    wire N__26989;
    wire N__26988;
    wire N__26983;
    wire N__26980;
    wire N__26977;
    wire N__26974;
    wire N__26971;
    wire N__26970;
    wire N__26969;
    wire N__26962;
    wire N__26961;
    wire N__26960;
    wire N__26957;
    wire N__26954;
    wire N__26951;
    wire N__26950;
    wire N__26947;
    wire N__26944;
    wire N__26939;
    wire N__26932;
    wire N__26929;
    wire N__26926;
    wire N__26923;
    wire N__26920;
    wire N__26919;
    wire N__26918;
    wire N__26915;
    wire N__26910;
    wire N__26907;
    wire N__26902;
    wire N__26899;
    wire N__26896;
    wire N__26893;
    wire N__26890;
    wire N__26887;
    wire N__26886;
    wire N__26883;
    wire N__26880;
    wire N__26877;
    wire N__26874;
    wire N__26873;
    wire N__26872;
    wire N__26871;
    wire N__26870;
    wire N__26867;
    wire N__26864;
    wire N__26861;
    wire N__26854;
    wire N__26851;
    wire N__26846;
    wire N__26839;
    wire N__26836;
    wire N__26833;
    wire N__26832;
    wire N__26831;
    wire N__26828;
    wire N__26825;
    wire N__26824;
    wire N__26821;
    wire N__26818;
    wire N__26815;
    wire N__26810;
    wire N__26807;
    wire N__26800;
    wire N__26797;
    wire N__26796;
    wire N__26795;
    wire N__26794;
    wire N__26791;
    wire N__26786;
    wire N__26785;
    wire N__26784;
    wire N__26781;
    wire N__26778;
    wire N__26775;
    wire N__26770;
    wire N__26761;
    wire N__26760;
    wire N__26757;
    wire N__26754;
    wire N__26749;
    wire N__26748;
    wire N__26745;
    wire N__26742;
    wire N__26739;
    wire N__26734;
    wire N__26733;
    wire N__26732;
    wire N__26731;
    wire N__26730;
    wire N__26729;
    wire N__26726;
    wire N__26719;
    wire N__26714;
    wire N__26713;
    wire N__26710;
    wire N__26705;
    wire N__26702;
    wire N__26699;
    wire N__26696;
    wire N__26693;
    wire N__26688;
    wire N__26685;
    wire N__26680;
    wire N__26679;
    wire N__26678;
    wire N__26677;
    wire N__26676;
    wire N__26675;
    wire N__26668;
    wire N__26667;
    wire N__26662;
    wire N__26659;
    wire N__26656;
    wire N__26653;
    wire N__26646;
    wire N__26641;
    wire N__26638;
    wire N__26637;
    wire N__26636;
    wire N__26631;
    wire N__26628;
    wire N__26623;
    wire N__26622;
    wire N__26621;
    wire N__26620;
    wire N__26611;
    wire N__26608;
    wire N__26605;
    wire N__26602;
    wire N__26599;
    wire N__26596;
    wire N__26593;
    wire N__26590;
    wire N__26587;
    wire N__26584;
    wire N__26583;
    wire N__26580;
    wire N__26577;
    wire N__26572;
    wire N__26569;
    wire N__26566;
    wire N__26565;
    wire N__26562;
    wire N__26559;
    wire N__26554;
    wire N__26551;
    wire N__26548;
    wire N__26545;
    wire N__26542;
    wire N__26541;
    wire N__26540;
    wire N__26537;
    wire N__26532;
    wire N__26527;
    wire N__26526;
    wire N__26523;
    wire N__26520;
    wire N__26515;
    wire N__26512;
    wire N__26511;
    wire N__26510;
    wire N__26509;
    wire N__26504;
    wire N__26503;
    wire N__26502;
    wire N__26501;
    wire N__26500;
    wire N__26497;
    wire N__26496;
    wire N__26495;
    wire N__26492;
    wire N__26491;
    wire N__26490;
    wire N__26487;
    wire N__26486;
    wire N__26483;
    wire N__26478;
    wire N__26469;
    wire N__26466;
    wire N__26461;
    wire N__26458;
    wire N__26455;
    wire N__26440;
    wire N__26439;
    wire N__26434;
    wire N__26431;
    wire N__26428;
    wire N__26427;
    wire N__26426;
    wire N__26425;
    wire N__26418;
    wire N__26417;
    wire N__26414;
    wire N__26411;
    wire N__26410;
    wire N__26409;
    wire N__26408;
    wire N__26407;
    wire N__26406;
    wire N__26403;
    wire N__26402;
    wire N__26401;
    wire N__26398;
    wire N__26395;
    wire N__26386;
    wire N__26383;
    wire N__26376;
    wire N__26365;
    wire N__26362;
    wire N__26359;
    wire N__26356;
    wire N__26355;
    wire N__26354;
    wire N__26351;
    wire N__26346;
    wire N__26341;
    wire N__26338;
    wire N__26337;
    wire N__26336;
    wire N__26335;
    wire N__26334;
    wire N__26333;
    wire N__26332;
    wire N__26331;
    wire N__26328;
    wire N__26321;
    wire N__26318;
    wire N__26317;
    wire N__26310;
    wire N__26305;
    wire N__26302;
    wire N__26301;
    wire N__26300;
    wire N__26299;
    wire N__26298;
    wire N__26297;
    wire N__26294;
    wire N__26293;
    wire N__26292;
    wire N__26289;
    wire N__26284;
    wire N__26273;
    wire N__26266;
    wire N__26257;
    wire N__26254;
    wire N__26251;
    wire N__26248;
    wire N__26245;
    wire N__26242;
    wire N__26239;
    wire N__26236;
    wire N__26233;
    wire N__26230;
    wire N__26229;
    wire N__26226;
    wire N__26225;
    wire N__26224;
    wire N__26223;
    wire N__26220;
    wire N__26217;
    wire N__26214;
    wire N__26209;
    wire N__26206;
    wire N__26197;
    wire N__26194;
    wire N__26193;
    wire N__26192;
    wire N__26189;
    wire N__26188;
    wire N__26185;
    wire N__26182;
    wire N__26179;
    wire N__26176;
    wire N__26171;
    wire N__26166;
    wire N__26161;
    wire N__26158;
    wire N__26157;
    wire N__26156;
    wire N__26153;
    wire N__26152;
    wire N__26151;
    wire N__26150;
    wire N__26149;
    wire N__26148;
    wire N__26147;
    wire N__26146;
    wire N__26145;
    wire N__26144;
    wire N__26143;
    wire N__26138;
    wire N__26135;
    wire N__26130;
    wire N__26127;
    wire N__26124;
    wire N__26121;
    wire N__26118;
    wire N__26115;
    wire N__26110;
    wire N__26107;
    wire N__26106;
    wire N__26105;
    wire N__26104;
    wire N__26103;
    wire N__26102;
    wire N__26101;
    wire N__26100;
    wire N__26099;
    wire N__26098;
    wire N__26097;
    wire N__26096;
    wire N__26095;
    wire N__26094;
    wire N__26093;
    wire N__26092;
    wire N__26091;
    wire N__26090;
    wire N__26089;
    wire N__26088;
    wire N__26087;
    wire N__26086;
    wire N__26085;
    wire N__26084;
    wire N__26083;
    wire N__26082;
    wire N__26081;
    wire N__26080;
    wire N__26079;
    wire N__26078;
    wire N__26077;
    wire N__26076;
    wire N__26075;
    wire N__26074;
    wire N__26073;
    wire N__26072;
    wire N__26071;
    wire N__26070;
    wire N__26069;
    wire N__26068;
    wire N__26067;
    wire N__26066;
    wire N__26065;
    wire N__26064;
    wire N__26063;
    wire N__26060;
    wire N__26057;
    wire N__26054;
    wire N__26051;
    wire N__26050;
    wire N__26049;
    wire N__26048;
    wire N__26047;
    wire N__26046;
    wire N__26045;
    wire N__26044;
    wire N__26043;
    wire N__26042;
    wire N__26041;
    wire N__26040;
    wire N__26039;
    wire N__26038;
    wire N__26037;
    wire N__26034;
    wire N__26031;
    wire N__26028;
    wire N__26025;
    wire N__26022;
    wire N__26019;
    wire N__25882;
    wire N__25879;
    wire N__25876;
    wire N__25875;
    wire N__25870;
    wire N__25867;
    wire N__25866;
    wire N__25865;
    wire N__25862;
    wire N__25857;
    wire N__25852;
    wire N__25851;
    wire N__25848;
    wire N__25845;
    wire N__25844;
    wire N__25843;
    wire N__25840;
    wire N__25837;
    wire N__25834;
    wire N__25831;
    wire N__25828;
    wire N__25823;
    wire N__25816;
    wire N__25813;
    wire N__25810;
    wire N__25809;
    wire N__25806;
    wire N__25803;
    wire N__25802;
    wire N__25799;
    wire N__25796;
    wire N__25793;
    wire N__25788;
    wire N__25783;
    wire N__25780;
    wire N__25779;
    wire N__25776;
    wire N__25775;
    wire N__25772;
    wire N__25769;
    wire N__25766;
    wire N__25763;
    wire N__25760;
    wire N__25753;
    wire N__25750;
    wire N__25747;
    wire N__25744;
    wire N__25741;
    wire N__25738;
    wire N__25735;
    wire N__25732;
    wire N__25729;
    wire N__25728;
    wire N__25725;
    wire N__25724;
    wire N__25721;
    wire N__25718;
    wire N__25715;
    wire N__25708;
    wire N__25705;
    wire N__25702;
    wire N__25699;
    wire N__25696;
    wire N__25693;
    wire N__25690;
    wire N__25687;
    wire N__25684;
    wire N__25683;
    wire N__25682;
    wire N__25677;
    wire N__25674;
    wire N__25671;
    wire N__25668;
    wire N__25665;
    wire N__25660;
    wire N__25659;
    wire N__25654;
    wire N__25651;
    wire N__25648;
    wire N__25645;
    wire N__25642;
    wire N__25639;
    wire N__25636;
    wire N__25633;
    wire N__25630;
    wire N__25629;
    wire N__25626;
    wire N__25625;
    wire N__25622;
    wire N__25619;
    wire N__25616;
    wire N__25609;
    wire N__25606;
    wire N__25603;
    wire N__25600;
    wire N__25597;
    wire N__25594;
    wire N__25591;
    wire N__25590;
    wire N__25587;
    wire N__25586;
    wire N__25583;
    wire N__25580;
    wire N__25577;
    wire N__25570;
    wire N__25567;
    wire N__25566;
    wire N__25565;
    wire N__25558;
    wire N__25555;
    wire N__25552;
    wire N__25551;
    wire N__25546;
    wire N__25543;
    wire N__25540;
    wire N__25537;
    wire N__25534;
    wire N__25533;
    wire N__25530;
    wire N__25527;
    wire N__25526;
    wire N__25523;
    wire N__25520;
    wire N__25517;
    wire N__25514;
    wire N__25511;
    wire N__25504;
    wire N__25501;
    wire N__25498;
    wire N__25495;
    wire N__25492;
    wire N__25491;
    wire N__25490;
    wire N__25489;
    wire N__25486;
    wire N__25479;
    wire N__25478;
    wire N__25477;
    wire N__25474;
    wire N__25471;
    wire N__25466;
    wire N__25461;
    wire N__25456;
    wire N__25453;
    wire N__25452;
    wire N__25447;
    wire N__25444;
    wire N__25441;
    wire N__25438;
    wire N__25435;
    wire N__25432;
    wire N__25429;
    wire N__25428;
    wire N__25427;
    wire N__25426;
    wire N__25425;
    wire N__25424;
    wire N__25423;
    wire N__25408;
    wire N__25405;
    wire N__25402;
    wire N__25399;
    wire N__25398;
    wire N__25397;
    wire N__25396;
    wire N__25395;
    wire N__25394;
    wire N__25391;
    wire N__25386;
    wire N__25381;
    wire N__25378;
    wire N__25377;
    wire N__25376;
    wire N__25375;
    wire N__25374;
    wire N__25373;
    wire N__25372;
    wire N__25363;
    wire N__25360;
    wire N__25357;
    wire N__25350;
    wire N__25347;
    wire N__25346;
    wire N__25345;
    wire N__25344;
    wire N__25341;
    wire N__25334;
    wire N__25331;
    wire N__25324;
    wire N__25315;
    wire N__25314;
    wire N__25313;
    wire N__25308;
    wire N__25305;
    wire N__25304;
    wire N__25303;
    wire N__25302;
    wire N__25301;
    wire N__25300;
    wire N__25297;
    wire N__25294;
    wire N__25291;
    wire N__25288;
    wire N__25283;
    wire N__25280;
    wire N__25279;
    wire N__25274;
    wire N__25273;
    wire N__25272;
    wire N__25269;
    wire N__25266;
    wire N__25261;
    wire N__25260;
    wire N__25257;
    wire N__25254;
    wire N__25251;
    wire N__25248;
    wire N__25241;
    wire N__25238;
    wire N__25225;
    wire N__25222;
    wire N__25219;
    wire N__25216;
    wire N__25213;
    wire N__25212;
    wire N__25211;
    wire N__25210;
    wire N__25201;
    wire N__25200;
    wire N__25199;
    wire N__25196;
    wire N__25193;
    wire N__25190;
    wire N__25185;
    wire N__25180;
    wire N__25179;
    wire N__25176;
    wire N__25173;
    wire N__25170;
    wire N__25167;
    wire N__25162;
    wire N__25161;
    wire N__25160;
    wire N__25157;
    wire N__25152;
    wire N__25147;
    wire N__25146;
    wire N__25143;
    wire N__25140;
    wire N__25137;
    wire N__25134;
    wire N__25133;
    wire N__25132;
    wire N__25131;
    wire N__25126;
    wire N__25119;
    wire N__25114;
    wire N__25111;
    wire N__25110;
    wire N__25109;
    wire N__25108;
    wire N__25105;
    wire N__25100;
    wire N__25097;
    wire N__25092;
    wire N__25089;
    wire N__25088;
    wire N__25085;
    wire N__25082;
    wire N__25079;
    wire N__25076;
    wire N__25069;
    wire N__25066;
    wire N__25063;
    wire N__25062;
    wire N__25061;
    wire N__25058;
    wire N__25053;
    wire N__25048;
    wire N__25047;
    wire N__25046;
    wire N__25045;
    wire N__25042;
    wire N__25041;
    wire N__25040;
    wire N__25039;
    wire N__25036;
    wire N__25033;
    wire N__25026;
    wire N__25025;
    wire N__25024;
    wire N__25023;
    wire N__25022;
    wire N__25021;
    wire N__25020;
    wire N__25019;
    wire N__25016;
    wire N__25013;
    wire N__25012;
    wire N__25011;
    wire N__25010;
    wire N__25009;
    wire N__25008;
    wire N__25005;
    wire N__25002;
    wire N__24999;
    wire N__24996;
    wire N__24987;
    wire N__24982;
    wire N__24979;
    wire N__24976;
    wire N__24973;
    wire N__24968;
    wire N__24965;
    wire N__24964;
    wire N__24961;
    wire N__24958;
    wire N__24953;
    wire N__24950;
    wire N__24947;
    wire N__24944;
    wire N__24935;
    wire N__24930;
    wire N__24927;
    wire N__24922;
    wire N__24919;
    wire N__24910;
    wire N__24901;
    wire N__24900;
    wire N__24899;
    wire N__24898;
    wire N__24897;
    wire N__24894;
    wire N__24891;
    wire N__24890;
    wire N__24889;
    wire N__24888;
    wire N__24887;
    wire N__24886;
    wire N__24885;
    wire N__24882;
    wire N__24879;
    wire N__24878;
    wire N__24875;
    wire N__24874;
    wire N__24871;
    wire N__24868;
    wire N__24865;
    wire N__24864;
    wire N__24863;
    wire N__24862;
    wire N__24861;
    wire N__24856;
    wire N__24849;
    wire N__24844;
    wire N__24841;
    wire N__24838;
    wire N__24835;
    wire N__24830;
    wire N__24827;
    wire N__24824;
    wire N__24819;
    wire N__24816;
    wire N__24815;
    wire N__24814;
    wire N__24813;
    wire N__24810;
    wire N__24807;
    wire N__24804;
    wire N__24803;
    wire N__24802;
    wire N__24797;
    wire N__24790;
    wire N__24787;
    wire N__24784;
    wire N__24779;
    wire N__24774;
    wire N__24767;
    wire N__24762;
    wire N__24757;
    wire N__24742;
    wire N__24739;
    wire N__24736;
    wire N__24733;
    wire N__24730;
    wire N__24727;
    wire N__24726;
    wire N__24725;
    wire N__24720;
    wire N__24717;
    wire N__24714;
    wire N__24711;
    wire N__24706;
    wire N__24705;
    wire N__24704;
    wire N__24703;
    wire N__24702;
    wire N__24699;
    wire N__24696;
    wire N__24695;
    wire N__24690;
    wire N__24689;
    wire N__24688;
    wire N__24687;
    wire N__24686;
    wire N__24685;
    wire N__24684;
    wire N__24683;
    wire N__24682;
    wire N__24681;
    wire N__24680;
    wire N__24679;
    wire N__24678;
    wire N__24677;
    wire N__24676;
    wire N__24675;
    wire N__24674;
    wire N__24673;
    wire N__24672;
    wire N__24671;
    wire N__24670;
    wire N__24669;
    wire N__24666;
    wire N__24663;
    wire N__24660;
    wire N__24657;
    wire N__24654;
    wire N__24651;
    wire N__24644;
    wire N__24637;
    wire N__24634;
    wire N__24631;
    wire N__24628;
    wire N__24627;
    wire N__24626;
    wire N__24623;
    wire N__24618;
    wire N__24615;
    wire N__24606;
    wire N__24599;
    wire N__24596;
    wire N__24591;
    wire N__24584;
    wire N__24579;
    wire N__24578;
    wire N__24577;
    wire N__24574;
    wire N__24569;
    wire N__24564;
    wire N__24557;
    wire N__24550;
    wire N__24547;
    wire N__24542;
    wire N__24537;
    wire N__24532;
    wire N__24525;
    wire N__24514;
    wire N__24513;
    wire N__24512;
    wire N__24509;
    wire N__24504;
    wire N__24499;
    wire N__24496;
    wire N__24495;
    wire N__24490;
    wire N__24487;
    wire N__24484;
    wire N__24481;
    wire N__24478;
    wire N__24477;
    wire N__24476;
    wire N__24475;
    wire N__24472;
    wire N__24469;
    wire N__24466;
    wire N__24463;
    wire N__24460;
    wire N__24457;
    wire N__24448;
    wire N__24447;
    wire N__24446;
    wire N__24445;
    wire N__24444;
    wire N__24443;
    wire N__24442;
    wire N__24441;
    wire N__24440;
    wire N__24437;
    wire N__24434;
    wire N__24429;
    wire N__24426;
    wire N__24423;
    wire N__24418;
    wire N__24417;
    wire N__24416;
    wire N__24415;
    wire N__24414;
    wire N__24411;
    wire N__24408;
    wire N__24401;
    wire N__24398;
    wire N__24395;
    wire N__24392;
    wire N__24387;
    wire N__24384;
    wire N__24379;
    wire N__24376;
    wire N__24371;
    wire N__24358;
    wire N__24357;
    wire N__24356;
    wire N__24351;
    wire N__24348;
    wire N__24347;
    wire N__24344;
    wire N__24341;
    wire N__24340;
    wire N__24337;
    wire N__24332;
    wire N__24329;
    wire N__24322;
    wire N__24321;
    wire N__24320;
    wire N__24317;
    wire N__24314;
    wire N__24311;
    wire N__24310;
    wire N__24309;
    wire N__24308;
    wire N__24301;
    wire N__24300;
    wire N__24297;
    wire N__24296;
    wire N__24295;
    wire N__24294;
    wire N__24291;
    wire N__24288;
    wire N__24285;
    wire N__24282;
    wire N__24275;
    wire N__24272;
    wire N__24271;
    wire N__24270;
    wire N__24267;
    wire N__24266;
    wire N__24263;
    wire N__24260;
    wire N__24255;
    wire N__24252;
    wire N__24247;
    wire N__24244;
    wire N__24241;
    wire N__24238;
    wire N__24235;
    wire N__24230;
    wire N__24217;
    wire N__24214;
    wire N__24211;
    wire N__24208;
    wire N__24207;
    wire N__24206;
    wire N__24203;
    wire N__24200;
    wire N__24197;
    wire N__24194;
    wire N__24191;
    wire N__24188;
    wire N__24185;
    wire N__24178;
    wire N__24177;
    wire N__24176;
    wire N__24173;
    wire N__24172;
    wire N__24169;
    wire N__24168;
    wire N__24165;
    wire N__24162;
    wire N__24159;
    wire N__24158;
    wire N__24157;
    wire N__24150;
    wire N__24145;
    wire N__24140;
    wire N__24133;
    wire N__24130;
    wire N__24127;
    wire N__24126;
    wire N__24123;
    wire N__24122;
    wire N__24121;
    wire N__24120;
    wire N__24113;
    wire N__24110;
    wire N__24107;
    wire N__24104;
    wire N__24101;
    wire N__24098;
    wire N__24095;
    wire N__24088;
    wire N__24085;
    wire N__24084;
    wire N__24081;
    wire N__24078;
    wire N__24073;
    wire N__24072;
    wire N__24069;
    wire N__24068;
    wire N__24061;
    wire N__24058;
    wire N__24057;
    wire N__24056;
    wire N__24055;
    wire N__24054;
    wire N__24053;
    wire N__24052;
    wire N__24047;
    wire N__24044;
    wire N__24035;
    wire N__24028;
    wire N__24025;
    wire N__24022;
    wire N__24019;
    wire N__24016;
    wire N__24013;
    wire N__24012;
    wire N__24011;
    wire N__24008;
    wire N__24007;
    wire N__24006;
    wire N__24005;
    wire N__24004;
    wire N__24003;
    wire N__24000;
    wire N__23997;
    wire N__23994;
    wire N__23991;
    wire N__23988;
    wire N__23985;
    wire N__23982;
    wire N__23977;
    wire N__23976;
    wire N__23973;
    wire N__23972;
    wire N__23969;
    wire N__23966;
    wire N__23963;
    wire N__23960;
    wire N__23955;
    wire N__23952;
    wire N__23949;
    wire N__23946;
    wire N__23937;
    wire N__23934;
    wire N__23923;
    wire N__23920;
    wire N__23917;
    wire N__23914;
    wire N__23913;
    wire N__23910;
    wire N__23907;
    wire N__23902;
    wire N__23899;
    wire N__23898;
    wire N__23895;
    wire N__23892;
    wire N__23889;
    wire N__23886;
    wire N__23883;
    wire N__23880;
    wire N__23877;
    wire N__23874;
    wire N__23869;
    wire N__23866;
    wire N__23863;
    wire N__23860;
    wire N__23857;
    wire N__23856;
    wire N__23855;
    wire N__23854;
    wire N__23851;
    wire N__23846;
    wire N__23843;
    wire N__23836;
    wire N__23833;
    wire N__23832;
    wire N__23831;
    wire N__23828;
    wire N__23827;
    wire N__23826;
    wire N__23825;
    wire N__23824;
    wire N__23819;
    wire N__23818;
    wire N__23817;
    wire N__23816;
    wire N__23815;
    wire N__23814;
    wire N__23813;
    wire N__23812;
    wire N__23807;
    wire N__23804;
    wire N__23799;
    wire N__23798;
    wire N__23795;
    wire N__23792;
    wire N__23789;
    wire N__23786;
    wire N__23785;
    wire N__23784;
    wire N__23781;
    wire N__23778;
    wire N__23777;
    wire N__23776;
    wire N__23775;
    wire N__23772;
    wire N__23769;
    wire N__23764;
    wire N__23761;
    wire N__23758;
    wire N__23749;
    wire N__23744;
    wire N__23741;
    wire N__23738;
    wire N__23731;
    wire N__23724;
    wire N__23721;
    wire N__23716;
    wire N__23709;
    wire N__23704;
    wire N__23699;
    wire N__23696;
    wire N__23693;
    wire N__23686;
    wire N__23685;
    wire N__23682;
    wire N__23679;
    wire N__23674;
    wire N__23671;
    wire N__23670;
    wire N__23665;
    wire N__23662;
    wire N__23659;
    wire N__23656;
    wire N__23655;
    wire N__23654;
    wire N__23647;
    wire N__23646;
    wire N__23645;
    wire N__23642;
    wire N__23639;
    wire N__23638;
    wire N__23637;
    wire N__23634;
    wire N__23631;
    wire N__23628;
    wire N__23623;
    wire N__23614;
    wire N__23611;
    wire N__23608;
    wire N__23605;
    wire N__23602;
    wire N__23599;
    wire N__23596;
    wire N__23595;
    wire N__23592;
    wire N__23589;
    wire N__23586;
    wire N__23581;
    wire N__23578;
    wire N__23575;
    wire N__23572;
    wire N__23571;
    wire N__23566;
    wire N__23563;
    wire N__23560;
    wire N__23557;
    wire N__23554;
    wire N__23551;
    wire N__23550;
    wire N__23549;
    wire N__23542;
    wire N__23539;
    wire N__23536;
    wire N__23533;
    wire N__23530;
    wire N__23527;
    wire N__23524;
    wire N__23521;
    wire N__23518;
    wire N__23515;
    wire N__23512;
    wire N__23509;
    wire N__23506;
    wire N__23503;
    wire N__23500;
    wire N__23497;
    wire N__23494;
    wire N__23491;
    wire N__23488;
    wire N__23485;
    wire N__23482;
    wire N__23479;
    wire N__23478;
    wire N__23477;
    wire N__23476;
    wire N__23473;
    wire N__23470;
    wire N__23465;
    wire N__23458;
    wire N__23457;
    wire N__23456;
    wire N__23455;
    wire N__23454;
    wire N__23453;
    wire N__23452;
    wire N__23449;
    wire N__23448;
    wire N__23447;
    wire N__23446;
    wire N__23445;
    wire N__23444;
    wire N__23441;
    wire N__23440;
    wire N__23439;
    wire N__23438;
    wire N__23437;
    wire N__23436;
    wire N__23435;
    wire N__23432;
    wire N__23431;
    wire N__23430;
    wire N__23423;
    wire N__23422;
    wire N__23415;
    wire N__23412;
    wire N__23405;
    wire N__23402;
    wire N__23397;
    wire N__23390;
    wire N__23389;
    wire N__23388;
    wire N__23385;
    wire N__23382;
    wire N__23381;
    wire N__23378;
    wire N__23377;
    wire N__23376;
    wire N__23375;
    wire N__23372;
    wire N__23369;
    wire N__23366;
    wire N__23363;
    wire N__23358;
    wire N__23351;
    wire N__23346;
    wire N__23345;
    wire N__23344;
    wire N__23343;
    wire N__23342;
    wire N__23341;
    wire N__23340;
    wire N__23337;
    wire N__23334;
    wire N__23331;
    wire N__23328;
    wire N__23327;
    wire N__23326;
    wire N__23321;
    wire N__23318;
    wire N__23315;
    wire N__23308;
    wire N__23301;
    wire N__23298;
    wire N__23295;
    wire N__23286;
    wire N__23277;
    wire N__23272;
    wire N__23261;
    wire N__23248;
    wire N__23247;
    wire N__23246;
    wire N__23241;
    wire N__23240;
    wire N__23239;
    wire N__23236;
    wire N__23235;
    wire N__23234;
    wire N__23233;
    wire N__23232;
    wire N__23229;
    wire N__23224;
    wire N__23223;
    wire N__23222;
    wire N__23221;
    wire N__23220;
    wire N__23217;
    wire N__23214;
    wire N__23207;
    wire N__23202;
    wire N__23199;
    wire N__23192;
    wire N__23187;
    wire N__23176;
    wire N__23175;
    wire N__23174;
    wire N__23171;
    wire N__23170;
    wire N__23163;
    wire N__23162;
    wire N__23161;
    wire N__23158;
    wire N__23157;
    wire N__23154;
    wire N__23147;
    wire N__23144;
    wire N__23141;
    wire N__23138;
    wire N__23131;
    wire N__23130;
    wire N__23127;
    wire N__23124;
    wire N__23121;
    wire N__23118;
    wire N__23113;
    wire N__23112;
    wire N__23109;
    wire N__23106;
    wire N__23105;
    wire N__23102;
    wire N__23097;
    wire N__23092;
    wire N__23091;
    wire N__23090;
    wire N__23087;
    wire N__23082;
    wire N__23077;
    wire N__23076;
    wire N__23075;
    wire N__23072;
    wire N__23069;
    wire N__23066;
    wire N__23059;
    wire N__23058;
    wire N__23057;
    wire N__23054;
    wire N__23051;
    wire N__23048;
    wire N__23045;
    wire N__23038;
    wire N__23037;
    wire N__23036;
    wire N__23033;
    wire N__23030;
    wire N__23027;
    wire N__23020;
    wire N__23019;
    wire N__23018;
    wire N__23015;
    wire N__23014;
    wire N__23011;
    wire N__23008;
    wire N__23003;
    wire N__22998;
    wire N__22995;
    wire N__22992;
    wire N__22989;
    wire N__22984;
    wire N__22983;
    wire N__22980;
    wire N__22979;
    wire N__22976;
    wire N__22973;
    wire N__22970;
    wire N__22963;
    wire N__22962;
    wire N__22961;
    wire N__22954;
    wire N__22953;
    wire N__22950;
    wire N__22947;
    wire N__22944;
    wire N__22941;
    wire N__22938;
    wire N__22935;
    wire N__22930;
    wire N__22929;
    wire N__22926;
    wire N__22925;
    wire N__22922;
    wire N__22919;
    wire N__22916;
    wire N__22909;
    wire N__22908;
    wire N__22907;
    wire N__22906;
    wire N__22897;
    wire N__22894;
    wire N__22891;
    wire N__22888;
    wire N__22885;
    wire N__22882;
    wire N__22881;
    wire N__22878;
    wire N__22875;
    wire N__22874;
    wire N__22873;
    wire N__22864;
    wire N__22861;
    wire N__22858;
    wire N__22855;
    wire N__22854;
    wire N__22851;
    wire N__22848;
    wire N__22843;
    wire N__22840;
    wire N__22837;
    wire N__22834;
    wire N__22831;
    wire N__22828;
    wire N__22827;
    wire N__22824;
    wire N__22821;
    wire N__22820;
    wire N__22815;
    wire N__22812;
    wire N__22807;
    wire N__22806;
    wire N__22803;
    wire N__22800;
    wire N__22797;
    wire N__22794;
    wire N__22793;
    wire N__22792;
    wire N__22787;
    wire N__22784;
    wire N__22781;
    wire N__22776;
    wire N__22773;
    wire N__22770;
    wire N__22765;
    wire N__22764;
    wire N__22761;
    wire N__22760;
    wire N__22757;
    wire N__22754;
    wire N__22751;
    wire N__22748;
    wire N__22745;
    wire N__22738;
    wire N__22735;
    wire N__22734;
    wire N__22733;
    wire N__22730;
    wire N__22727;
    wire N__22724;
    wire N__22721;
    wire N__22714;
    wire N__22713;
    wire N__22712;
    wire N__22711;
    wire N__22702;
    wire N__22699;
    wire N__22696;
    wire N__22693;
    wire N__22690;
    wire N__22689;
    wire N__22688;
    wire N__22685;
    wire N__22682;
    wire N__22679;
    wire N__22676;
    wire N__22669;
    wire N__22666;
    wire N__22665;
    wire N__22662;
    wire N__22661;
    wire N__22658;
    wire N__22655;
    wire N__22652;
    wire N__22649;
    wire N__22642;
    wire N__22639;
    wire N__22636;
    wire N__22633;
    wire N__22632;
    wire N__22631;
    wire N__22628;
    wire N__22623;
    wire N__22618;
    wire N__22615;
    wire N__22614;
    wire N__22613;
    wire N__22610;
    wire N__22605;
    wire N__22600;
    wire N__22597;
    wire N__22596;
    wire N__22595;
    wire N__22594;
    wire N__22593;
    wire N__22582;
    wire N__22579;
    wire N__22578;
    wire N__22577;
    wire N__22576;
    wire N__22569;
    wire N__22566;
    wire N__22561;
    wire N__22560;
    wire N__22557;
    wire N__22556;
    wire N__22551;
    wire N__22548;
    wire N__22543;
    wire N__22540;
    wire N__22539;
    wire N__22538;
    wire N__22537;
    wire N__22534;
    wire N__22525;
    wire N__22522;
    wire N__22521;
    wire N__22520;
    wire N__22519;
    wire N__22516;
    wire N__22515;
    wire N__22506;
    wire N__22503;
    wire N__22498;
    wire N__22495;
    wire N__22492;
    wire N__22489;
    wire N__22488;
    wire N__22487;
    wire N__22486;
    wire N__22481;
    wire N__22478;
    wire N__22475;
    wire N__22472;
    wire N__22469;
    wire N__22462;
    wire N__22461;
    wire N__22460;
    wire N__22459;
    wire N__22456;
    wire N__22455;
    wire N__22450;
    wire N__22447;
    wire N__22442;
    wire N__22439;
    wire N__22436;
    wire N__22429;
    wire N__22428;
    wire N__22427;
    wire N__22426;
    wire N__22425;
    wire N__22424;
    wire N__22423;
    wire N__22416;
    wire N__22409;
    wire N__22406;
    wire N__22399;
    wire N__22398;
    wire N__22397;
    wire N__22396;
    wire N__22395;
    wire N__22390;
    wire N__22383;
    wire N__22378;
    wire N__22375;
    wire N__22374;
    wire N__22371;
    wire N__22370;
    wire N__22367;
    wire N__22364;
    wire N__22359;
    wire N__22354;
    wire N__22353;
    wire N__22352;
    wire N__22351;
    wire N__22350;
    wire N__22343;
    wire N__22340;
    wire N__22337;
    wire N__22332;
    wire N__22327;
    wire N__22326;
    wire N__22323;
    wire N__22322;
    wire N__22319;
    wire N__22316;
    wire N__22313;
    wire N__22312;
    wire N__22307;
    wire N__22304;
    wire N__22301;
    wire N__22294;
    wire N__22293;
    wire N__22292;
    wire N__22285;
    wire N__22282;
    wire N__22281;
    wire N__22280;
    wire N__22277;
    wire N__22272;
    wire N__22269;
    wire N__22264;
    wire N__22261;
    wire N__22260;
    wire N__22259;
    wire N__22256;
    wire N__22251;
    wire N__22248;
    wire N__22243;
    wire N__22242;
    wire N__22241;
    wire N__22236;
    wire N__22235;
    wire N__22232;
    wire N__22229;
    wire N__22226;
    wire N__22219;
    wire N__22216;
    wire N__22215;
    wire N__22214;
    wire N__22213;
    wire N__22208;
    wire N__22205;
    wire N__22202;
    wire N__22195;
    wire N__22194;
    wire N__22193;
    wire N__22192;
    wire N__22187;
    wire N__22184;
    wire N__22181;
    wire N__22174;
    wire N__22173;
    wire N__22172;
    wire N__22171;
    wire N__22170;
    wire N__22159;
    wire N__22156;
    wire N__22153;
    wire N__22150;
    wire N__22147;
    wire N__22146;
    wire N__22143;
    wire N__22140;
    wire N__22135;
    wire N__22132;
    wire N__22129;
    wire N__22128;
    wire N__22127;
    wire N__22124;
    wire N__22121;
    wire N__22118;
    wire N__22111;
    wire N__22110;
    wire N__22109;
    wire N__22106;
    wire N__22103;
    wire N__22096;
    wire N__22093;
    wire N__22092;
    wire N__22091;
    wire N__22090;
    wire N__22083;
    wire N__22080;
    wire N__22075;
    wire N__22072;
    wire N__22071;
    wire N__22068;
    wire N__22065;
    wire N__22062;
    wire N__22057;
    wire N__22056;
    wire N__22055;
    wire N__22052;
    wire N__22049;
    wire N__22046;
    wire N__22039;
    wire N__22036;
    wire N__22035;
    wire N__22034;
    wire N__22033;
    wire N__22026;
    wire N__22023;
    wire N__22018;
    wire N__22015;
    wire N__22012;
    wire N__22009;
    wire N__22006;
    wire N__22003;
    wire N__22000;
    wire N__21999;
    wire N__21996;
    wire N__21995;
    wire N__21992;
    wire N__21991;
    wire N__21988;
    wire N__21987;
    wire N__21986;
    wire N__21983;
    wire N__21980;
    wire N__21977;
    wire N__21974;
    wire N__21971;
    wire N__21966;
    wire N__21963;
    wire N__21960;
    wire N__21957;
    wire N__21954;
    wire N__21949;
    wire N__21946;
    wire N__21937;
    wire N__21936;
    wire N__21935;
    wire N__21932;
    wire N__21929;
    wire N__21926;
    wire N__21925;
    wire N__21924;
    wire N__21919;
    wire N__21918;
    wire N__21915;
    wire N__21910;
    wire N__21907;
    wire N__21904;
    wire N__21895;
    wire N__21892;
    wire N__21891;
    wire N__21888;
    wire N__21885;
    wire N__21882;
    wire N__21877;
    wire N__21876;
    wire N__21873;
    wire N__21872;
    wire N__21871;
    wire N__21868;
    wire N__21865;
    wire N__21862;
    wire N__21859;
    wire N__21852;
    wire N__21849;
    wire N__21846;
    wire N__21841;
    wire N__21838;
    wire N__21837;
    wire N__21834;
    wire N__21833;
    wire N__21832;
    wire N__21831;
    wire N__21828;
    wire N__21825;
    wire N__21820;
    wire N__21819;
    wire N__21816;
    wire N__21813;
    wire N__21810;
    wire N__21807;
    wire N__21802;
    wire N__21793;
    wire N__21790;
    wire N__21787;
    wire N__21784;
    wire N__21781;
    wire N__21780;
    wire N__21777;
    wire N__21774;
    wire N__21771;
    wire N__21768;
    wire N__21767;
    wire N__21766;
    wire N__21765;
    wire N__21764;
    wire N__21763;
    wire N__21760;
    wire N__21757;
    wire N__21756;
    wire N__21753;
    wire N__21750;
    wire N__21749;
    wire N__21742;
    wire N__21739;
    wire N__21736;
    wire N__21727;
    wire N__21718;
    wire N__21715;
    wire N__21712;
    wire N__21709;
    wire N__21706;
    wire N__21703;
    wire N__21700;
    wire N__21699;
    wire N__21698;
    wire N__21697;
    wire N__21696;
    wire N__21695;
    wire N__21692;
    wire N__21689;
    wire N__21686;
    wire N__21685;
    wire N__21684;
    wire N__21683;
    wire N__21680;
    wire N__21675;
    wire N__21672;
    wire N__21669;
    wire N__21660;
    wire N__21649;
    wire N__21646;
    wire N__21643;
    wire N__21640;
    wire N__21637;
    wire N__21634;
    wire N__21631;
    wire N__21628;
    wire N__21625;
    wire N__21624;
    wire N__21623;
    wire N__21622;
    wire N__21621;
    wire N__21620;
    wire N__21619;
    wire N__21618;
    wire N__21617;
    wire N__21616;
    wire N__21615;
    wire N__21614;
    wire N__21611;
    wire N__21610;
    wire N__21609;
    wire N__21608;
    wire N__21607;
    wire N__21606;
    wire N__21603;
    wire N__21598;
    wire N__21581;
    wire N__21578;
    wire N__21577;
    wire N__21576;
    wire N__21575;
    wire N__21574;
    wire N__21573;
    wire N__21572;
    wire N__21569;
    wire N__21568;
    wire N__21565;
    wire N__21562;
    wire N__21559;
    wire N__21556;
    wire N__21553;
    wire N__21550;
    wire N__21547;
    wire N__21544;
    wire N__21537;
    wire N__21536;
    wire N__21529;
    wire N__21522;
    wire N__21521;
    wire N__21520;
    wire N__21519;
    wire N__21518;
    wire N__21517;
    wire N__21516;
    wire N__21515;
    wire N__21514;
    wire N__21513;
    wire N__21508;
    wire N__21501;
    wire N__21496;
    wire N__21493;
    wire N__21490;
    wire N__21485;
    wire N__21470;
    wire N__21465;
    wire N__21462;
    wire N__21445;
    wire N__21444;
    wire N__21443;
    wire N__21442;
    wire N__21441;
    wire N__21438;
    wire N__21435;
    wire N__21430;
    wire N__21427;
    wire N__21420;
    wire N__21415;
    wire N__21414;
    wire N__21411;
    wire N__21408;
    wire N__21407;
    wire N__21406;
    wire N__21403;
    wire N__21400;
    wire N__21395;
    wire N__21394;
    wire N__21393;
    wire N__21392;
    wire N__21391;
    wire N__21390;
    wire N__21389;
    wire N__21384;
    wire N__21381;
    wire N__21376;
    wire N__21367;
    wire N__21358;
    wire N__21355;
    wire N__21352;
    wire N__21351;
    wire N__21348;
    wire N__21347;
    wire N__21346;
    wire N__21343;
    wire N__21340;
    wire N__21335;
    wire N__21330;
    wire N__21325;
    wire N__21322;
    wire N__21319;
    wire N__21316;
    wire N__21313;
    wire N__21310;
    wire N__21307;
    wire N__21304;
    wire N__21301;
    wire N__21298;
    wire N__21295;
    wire N__21292;
    wire N__21291;
    wire N__21290;
    wire N__21287;
    wire N__21286;
    wire N__21281;
    wire N__21278;
    wire N__21275;
    wire N__21268;
    wire N__21267;
    wire N__21266;
    wire N__21265;
    wire N__21264;
    wire N__21261;
    wire N__21260;
    wire N__21259;
    wire N__21254;
    wire N__21251;
    wire N__21250;
    wire N__21247;
    wire N__21246;
    wire N__21245;
    wire N__21244;
    wire N__21241;
    wire N__21238;
    wire N__21235;
    wire N__21234;
    wire N__21231;
    wire N__21228;
    wire N__21223;
    wire N__21222;
    wire N__21219;
    wire N__21218;
    wire N__21215;
    wire N__21212;
    wire N__21207;
    wire N__21204;
    wire N__21201;
    wire N__21194;
    wire N__21191;
    wire N__21188;
    wire N__21185;
    wire N__21182;
    wire N__21179;
    wire N__21176;
    wire N__21171;
    wire N__21168;
    wire N__21165;
    wire N__21160;
    wire N__21157;
    wire N__21152;
    wire N__21147;
    wire N__21136;
    wire N__21133;
    wire N__21130;
    wire N__21127;
    wire N__21124;
    wire N__21121;
    wire N__21118;
    wire N__21115;
    wire N__21112;
    wire N__21111;
    wire N__21110;
    wire N__21109;
    wire N__21108;
    wire N__21107;
    wire N__21104;
    wire N__21099;
    wire N__21098;
    wire N__21097;
    wire N__21096;
    wire N__21095;
    wire N__21094;
    wire N__21093;
    wire N__21092;
    wire N__21091;
    wire N__21090;
    wire N__21087;
    wire N__21084;
    wire N__21081;
    wire N__21076;
    wire N__21073;
    wire N__21072;
    wire N__21071;
    wire N__21054;
    wire N__21051;
    wire N__21048;
    wire N__21045;
    wire N__21044;
    wire N__21043;
    wire N__21042;
    wire N__21041;
    wire N__21040;
    wire N__21039;
    wire N__21038;
    wire N__21037;
    wire N__21036;
    wire N__21035;
    wire N__21034;
    wire N__21033;
    wire N__21032;
    wire N__21031;
    wire N__21030;
    wire N__21029;
    wire N__21028;
    wire N__21023;
    wire N__21020;
    wire N__21017;
    wire N__21008;
    wire N__21001;
    wire N__20990;
    wire N__20985;
    wire N__20970;
    wire N__20967;
    wire N__20950;
    wire N__20949;
    wire N__20946;
    wire N__20941;
    wire N__20940;
    wire N__20939;
    wire N__20938;
    wire N__20937;
    wire N__20936;
    wire N__20935;
    wire N__20932;
    wire N__20929;
    wire N__20926;
    wire N__20923;
    wire N__20916;
    wire N__20913;
    wire N__20910;
    wire N__20907;
    wire N__20904;
    wire N__20901;
    wire N__20900;
    wire N__20895;
    wire N__20892;
    wire N__20891;
    wire N__20886;
    wire N__20883;
    wire N__20880;
    wire N__20877;
    wire N__20874;
    wire N__20871;
    wire N__20860;
    wire N__20857;
    wire N__20854;
    wire N__20851;
    wire N__20848;
    wire N__20845;
    wire N__20842;
    wire N__20839;
    wire N__20838;
    wire N__20835;
    wire N__20832;
    wire N__20829;
    wire N__20824;
    wire N__20821;
    wire N__20818;
    wire N__20815;
    wire N__20814;
    wire N__20813;
    wire N__20812;
    wire N__20811;
    wire N__20810;
    wire N__20809;
    wire N__20808;
    wire N__20807;
    wire N__20806;
    wire N__20805;
    wire N__20802;
    wire N__20799;
    wire N__20796;
    wire N__20795;
    wire N__20794;
    wire N__20793;
    wire N__20792;
    wire N__20789;
    wire N__20786;
    wire N__20783;
    wire N__20780;
    wire N__20777;
    wire N__20774;
    wire N__20771;
    wire N__20768;
    wire N__20767;
    wire N__20764;
    wire N__20761;
    wire N__20758;
    wire N__20757;
    wire N__20756;
    wire N__20755;
    wire N__20752;
    wire N__20751;
    wire N__20748;
    wire N__20747;
    wire N__20746;
    wire N__20743;
    wire N__20742;
    wire N__20739;
    wire N__20730;
    wire N__20721;
    wire N__20718;
    wire N__20713;
    wire N__20710;
    wire N__20705;
    wire N__20698;
    wire N__20685;
    wire N__20668;
    wire N__20667;
    wire N__20666;
    wire N__20665;
    wire N__20664;
    wire N__20663;
    wire N__20662;
    wire N__20661;
    wire N__20660;
    wire N__20659;
    wire N__20658;
    wire N__20657;
    wire N__20654;
    wire N__20653;
    wire N__20644;
    wire N__20635;
    wire N__20634;
    wire N__20631;
    wire N__20628;
    wire N__20627;
    wire N__20624;
    wire N__20623;
    wire N__20622;
    wire N__20619;
    wire N__20616;
    wire N__20611;
    wire N__20598;
    wire N__20595;
    wire N__20592;
    wire N__20585;
    wire N__20578;
    wire N__20575;
    wire N__20572;
    wire N__20569;
    wire N__20566;
    wire N__20563;
    wire N__20562;
    wire N__20561;
    wire N__20560;
    wire N__20557;
    wire N__20554;
    wire N__20551;
    wire N__20548;
    wire N__20539;
    wire N__20536;
    wire N__20533;
    wire N__20530;
    wire N__20529;
    wire N__20524;
    wire N__20521;
    wire N__20518;
    wire N__20517;
    wire N__20516;
    wire N__20515;
    wire N__20508;
    wire N__20507;
    wire N__20506;
    wire N__20503;
    wire N__20500;
    wire N__20495;
    wire N__20492;
    wire N__20487;
    wire N__20484;
    wire N__20481;
    wire N__20476;
    wire N__20475;
    wire N__20472;
    wire N__20469;
    wire N__20466;
    wire N__20463;
    wire N__20458;
    wire N__20457;
    wire N__20454;
    wire N__20451;
    wire N__20448;
    wire N__20445;
    wire N__20442;
    wire N__20437;
    wire N__20434;
    wire N__20433;
    wire N__20428;
    wire N__20425;
    wire N__20424;
    wire N__20423;
    wire N__20422;
    wire N__20419;
    wire N__20412;
    wire N__20409;
    wire N__20406;
    wire N__20401;
    wire N__20398;
    wire N__20397;
    wire N__20396;
    wire N__20395;
    wire N__20394;
    wire N__20393;
    wire N__20392;
    wire N__20389;
    wire N__20388;
    wire N__20385;
    wire N__20382;
    wire N__20379;
    wire N__20374;
    wire N__20371;
    wire N__20370;
    wire N__20369;
    wire N__20362;
    wire N__20361;
    wire N__20360;
    wire N__20357;
    wire N__20352;
    wire N__20349;
    wire N__20346;
    wire N__20343;
    wire N__20340;
    wire N__20335;
    wire N__20334;
    wire N__20329;
    wire N__20324;
    wire N__20321;
    wire N__20316;
    wire N__20313;
    wire N__20308;
    wire N__20299;
    wire N__20296;
    wire N__20295;
    wire N__20292;
    wire N__20289;
    wire N__20284;
    wire N__20283;
    wire N__20280;
    wire N__20277;
    wire N__20274;
    wire N__20271;
    wire N__20268;
    wire N__20263;
    wire N__20260;
    wire N__20257;
    wire N__20254;
    wire N__20251;
    wire N__20248;
    wire N__20245;
    wire N__20242;
    wire N__20239;
    wire N__20236;
    wire N__20235;
    wire N__20230;
    wire N__20227;
    wire N__20224;
    wire N__20223;
    wire N__20220;
    wire N__20217;
    wire N__20212;
    wire N__20209;
    wire N__20206;
    wire N__20203;
    wire N__20200;
    wire N__20197;
    wire N__20194;
    wire N__20191;
    wire N__20188;
    wire N__20185;
    wire N__20182;
    wire N__20179;
    wire N__20178;
    wire N__20173;
    wire N__20170;
    wire N__20169;
    wire N__20168;
    wire N__20167;
    wire N__20166;
    wire N__20165;
    wire N__20164;
    wire N__20161;
    wire N__20154;
    wire N__20147;
    wire N__20144;
    wire N__20141;
    wire N__20138;
    wire N__20135;
    wire N__20130;
    wire N__20125;
    wire N__20122;
    wire N__20119;
    wire N__20118;
    wire N__20115;
    wire N__20112;
    wire N__20107;
    wire N__20106;
    wire N__20103;
    wire N__20100;
    wire N__20095;
    wire N__20092;
    wire N__20089;
    wire N__20086;
    wire N__20083;
    wire N__20080;
    wire N__20077;
    wire N__20076;
    wire N__20075;
    wire N__20074;
    wire N__20073;
    wire N__20072;
    wire N__20071;
    wire N__20062;
    wire N__20055;
    wire N__20052;
    wire N__20047;
    wire N__20046;
    wire N__20045;
    wire N__20044;
    wire N__20043;
    wire N__20042;
    wire N__20041;
    wire N__20040;
    wire N__20031;
    wire N__20030;
    wire N__20021;
    wire N__20018;
    wire N__20015;
    wire N__20008;
    wire N__20007;
    wire N__20006;
    wire N__20005;
    wire N__20002;
    wire N__19993;
    wire N__19992;
    wire N__19991;
    wire N__19988;
    wire N__19987;
    wire N__19984;
    wire N__19983;
    wire N__19980;
    wire N__19979;
    wire N__19976;
    wire N__19973;
    wire N__19966;
    wire N__19963;
    wire N__19954;
    wire N__19951;
    wire N__19950;
    wire N__19949;
    wire N__19948;
    wire N__19945;
    wire N__19942;
    wire N__19939;
    wire N__19938;
    wire N__19937;
    wire N__19934;
    wire N__19933;
    wire N__19924;
    wire N__19923;
    wire N__19916;
    wire N__19913;
    wire N__19910;
    wire N__19903;
    wire N__19900;
    wire N__19897;
    wire N__19896;
    wire N__19895;
    wire N__19894;
    wire N__19893;
    wire N__19890;
    wire N__19889;
    wire N__19888;
    wire N__19887;
    wire N__19886;
    wire N__19885;
    wire N__19884;
    wire N__19883;
    wire N__19882;
    wire N__19881;
    wire N__19880;
    wire N__19879;
    wire N__19878;
    wire N__19877;
    wire N__19876;
    wire N__19875;
    wire N__19870;
    wire N__19865;
    wire N__19858;
    wire N__19857;
    wire N__19856;
    wire N__19855;
    wire N__19852;
    wire N__19851;
    wire N__19850;
    wire N__19849;
    wire N__19848;
    wire N__19845;
    wire N__19840;
    wire N__19835;
    wire N__19828;
    wire N__19821;
    wire N__19820;
    wire N__19817;
    wire N__19810;
    wire N__19807;
    wire N__19802;
    wire N__19797;
    wire N__19790;
    wire N__19783;
    wire N__19778;
    wire N__19773;
    wire N__19770;
    wire N__19761;
    wire N__19758;
    wire N__19755;
    wire N__19750;
    wire N__19741;
    wire N__19740;
    wire N__19739;
    wire N__19738;
    wire N__19737;
    wire N__19736;
    wire N__19733;
    wire N__19730;
    wire N__19727;
    wire N__19726;
    wire N__19723;
    wire N__19722;
    wire N__19713;
    wire N__19704;
    wire N__19699;
    wire N__19696;
    wire N__19695;
    wire N__19690;
    wire N__19687;
    wire N__19684;
    wire N__19683;
    wire N__19682;
    wire N__19681;
    wire N__19672;
    wire N__19671;
    wire N__19670;
    wire N__19669;
    wire N__19668;
    wire N__19667;
    wire N__19666;
    wire N__19665;
    wire N__19664;
    wire N__19661;
    wire N__19660;
    wire N__19659;
    wire N__19646;
    wire N__19645;
    wire N__19644;
    wire N__19639;
    wire N__19636;
    wire N__19631;
    wire N__19628;
    wire N__19623;
    wire N__19612;
    wire N__19609;
    wire N__19608;
    wire N__19605;
    wire N__19604;
    wire N__19603;
    wire N__19594;
    wire N__19591;
    wire N__19590;
    wire N__19589;
    wire N__19588;
    wire N__19587;
    wire N__19584;
    wire N__19581;
    wire N__19576;
    wire N__19573;
    wire N__19564;
    wire N__19563;
    wire N__19562;
    wire N__19561;
    wire N__19560;
    wire N__19559;
    wire N__19556;
    wire N__19549;
    wire N__19544;
    wire N__19543;
    wire N__19536;
    wire N__19533;
    wire N__19530;
    wire N__19527;
    wire N__19522;
    wire N__19519;
    wire N__19516;
    wire N__19513;
    wire N__19510;
    wire N__19507;
    wire N__19504;
    wire N__19501;
    wire N__19498;
    wire N__19497;
    wire N__19496;
    wire N__19495;
    wire N__19494;
    wire N__19493;
    wire N__19492;
    wire N__19491;
    wire N__19488;
    wire N__19487;
    wire N__19484;
    wire N__19483;
    wire N__19480;
    wire N__19477;
    wire N__19474;
    wire N__19473;
    wire N__19468;
    wire N__19465;
    wire N__19460;
    wire N__19459;
    wire N__19458;
    wire N__19453;
    wire N__19448;
    wire N__19445;
    wire N__19442;
    wire N__19439;
    wire N__19438;
    wire N__19437;
    wire N__19436;
    wire N__19435;
    wire N__19432;
    wire N__19429;
    wire N__19426;
    wire N__19425;
    wire N__19422;
    wire N__19415;
    wire N__19410;
    wire N__19407;
    wire N__19402;
    wire N__19399;
    wire N__19394;
    wire N__19391;
    wire N__19386;
    wire N__19369;
    wire N__19366;
    wire N__19363;
    wire N__19360;
    wire N__19359;
    wire N__19358;
    wire N__19357;
    wire N__19356;
    wire N__19355;
    wire N__19354;
    wire N__19353;
    wire N__19344;
    wire N__19335;
    wire N__19330;
    wire N__19327;
    wire N__19324;
    wire N__19321;
    wire N__19318;
    wire N__19317;
    wire N__19316;
    wire N__19315;
    wire N__19312;
    wire N__19311;
    wire N__19310;
    wire N__19307;
    wire N__19306;
    wire N__19305;
    wire N__19304;
    wire N__19301;
    wire N__19298;
    wire N__19289;
    wire N__19286;
    wire N__19277;
    wire N__19270;
    wire N__19269;
    wire N__19268;
    wire N__19267;
    wire N__19266;
    wire N__19265;
    wire N__19264;
    wire N__19263;
    wire N__19254;
    wire N__19245;
    wire N__19240;
    wire N__19239;
    wire N__19238;
    wire N__19231;
    wire N__19228;
    wire N__19227;
    wire N__19226;
    wire N__19219;
    wire N__19218;
    wire N__19215;
    wire N__19212;
    wire N__19209;
    wire N__19204;
    wire N__19201;
    wire N__19198;
    wire N__19195;
    wire N__19192;
    wire N__19191;
    wire N__19188;
    wire N__19187;
    wire N__19186;
    wire N__19183;
    wire N__19176;
    wire N__19173;
    wire N__19172;
    wire N__19171;
    wire N__19168;
    wire N__19165;
    wire N__19162;
    wire N__19159;
    wire N__19154;
    wire N__19147;
    wire N__19144;
    wire N__19141;
    wire N__19140;
    wire N__19139;
    wire N__19136;
    wire N__19131;
    wire N__19128;
    wire N__19123;
    wire N__19120;
    wire N__19117;
    wire N__19114;
    wire N__19111;
    wire N__19108;
    wire N__19105;
    wire N__19102;
    wire N__19099;
    wire N__19096;
    wire N__19093;
    wire N__19090;
    wire N__19087;
    wire N__19084;
    wire N__19081;
    wire N__19078;
    wire N__19075;
    wire N__19072;
    wire N__19069;
    wire N__19068;
    wire N__19065;
    wire N__19064;
    wire N__19063;
    wire N__19062;
    wire N__19051;
    wire N__19050;
    wire N__19049;
    wire N__19046;
    wire N__19041;
    wire N__19036;
    wire N__19035;
    wire N__19034;
    wire N__19031;
    wire N__19030;
    wire N__19027;
    wire N__19024;
    wire N__19023;
    wire N__19018;
    wire N__19015;
    wire N__19010;
    wire N__19007;
    wire N__19004;
    wire N__18997;
    wire N__18994;
    wire N__18993;
    wire N__18992;
    wire N__18991;
    wire N__18988;
    wire N__18983;
    wire N__18980;
    wire N__18973;
    wire N__18970;
    wire N__18969;
    wire N__18968;
    wire N__18967;
    wire N__18964;
    wire N__18963;
    wire N__18962;
    wire N__18955;
    wire N__18952;
    wire N__18947;
    wire N__18940;
    wire N__18937;
    wire N__18934;
    wire N__18933;
    wire N__18930;
    wire N__18927;
    wire N__18924;
    wire N__18919;
    wire N__18918;
    wire N__18915;
    wire N__18912;
    wire N__18909;
    wire N__18906;
    wire N__18903;
    wire N__18898;
    wire N__18895;
    wire N__18892;
    wire N__18891;
    wire N__18888;
    wire N__18883;
    wire N__18880;
    wire N__18879;
    wire N__18878;
    wire N__18871;
    wire N__18868;
    wire N__18865;
    wire N__18864;
    wire N__18863;
    wire N__18858;
    wire N__18855;
    wire N__18852;
    wire N__18847;
    wire N__18844;
    wire N__18841;
    wire N__18838;
    wire N__18835;
    wire N__18832;
    wire N__18829;
    wire N__18826;
    wire N__18823;
    wire N__18820;
    wire N__18817;
    wire N__18814;
    wire N__18811;
    wire N__18808;
    wire N__18805;
    wire N__18802;
    wire N__18801;
    wire N__18800;
    wire N__18799;
    wire N__18798;
    wire N__18787;
    wire N__18786;
    wire N__18785;
    wire N__18782;
    wire N__18779;
    wire N__18776;
    wire N__18775;
    wire N__18774;
    wire N__18773;
    wire N__18772;
    wire N__18771;
    wire N__18764;
    wire N__18761;
    wire N__18752;
    wire N__18751;
    wire N__18750;
    wire N__18749;
    wire N__18748;
    wire N__18745;
    wire N__18742;
    wire N__18739;
    wire N__18734;
    wire N__18731;
    wire N__18728;
    wire N__18715;
    wire N__18712;
    wire N__18709;
    wire N__18706;
    wire N__18703;
    wire N__18700;
    wire N__18697;
    wire N__18694;
    wire N__18691;
    wire N__18690;
    wire N__18689;
    wire N__18688;
    wire N__18685;
    wire N__18678;
    wire N__18673;
    wire N__18672;
    wire N__18671;
    wire N__18670;
    wire N__18667;
    wire N__18664;
    wire N__18661;
    wire N__18656;
    wire N__18651;
    wire N__18646;
    wire N__18645;
    wire N__18644;
    wire N__18643;
    wire N__18640;
    wire N__18633;
    wire N__18628;
    wire N__18625;
    wire N__18622;
    wire N__18621;
    wire N__18620;
    wire N__18613;
    wire N__18610;
    wire N__18609;
    wire N__18608;
    wire N__18605;
    wire N__18604;
    wire N__18603;
    wire N__18602;
    wire N__18601;
    wire N__18598;
    wire N__18595;
    wire N__18594;
    wire N__18593;
    wire N__18592;
    wire N__18585;
    wire N__18582;
    wire N__18577;
    wire N__18568;
    wire N__18559;
    wire N__18558;
    wire N__18557;
    wire N__18556;
    wire N__18555;
    wire N__18554;
    wire N__18547;
    wire N__18540;
    wire N__18535;
    wire N__18532;
    wire N__18529;
    wire N__18526;
    wire N__18523;
    wire N__18520;
    wire N__18517;
    wire N__18514;
    wire N__18513;
    wire N__18508;
    wire N__18505;
    wire N__18502;
    wire N__18501;
    wire N__18500;
    wire N__18495;
    wire N__18492;
    wire N__18487;
    wire N__18486;
    wire N__18483;
    wire N__18480;
    wire N__18479;
    wire N__18476;
    wire N__18471;
    wire N__18468;
    wire N__18463;
    wire N__18460;
    wire N__18457;
    wire N__18454;
    wire N__18453;
    wire N__18452;
    wire N__18451;
    wire N__18450;
    wire N__18447;
    wire N__18440;
    wire N__18437;
    wire N__18430;
    wire N__18429;
    wire N__18428;
    wire N__18427;
    wire N__18424;
    wire N__18421;
    wire N__18416;
    wire N__18409;
    wire N__18406;
    wire N__18403;
    wire N__18400;
    wire N__18397;
    wire N__18394;
    wire N__18391;
    wire N__18388;
    wire N__18385;
    wire N__18382;
    wire N__18379;
    wire N__18376;
    wire N__18375;
    wire N__18372;
    wire N__18371;
    wire N__18368;
    wire N__18367;
    wire N__18366;
    wire N__18361;
    wire N__18358;
    wire N__18353;
    wire N__18348;
    wire N__18343;
    wire N__18340;
    wire N__18337;
    wire N__18334;
    wire N__18331;
    wire N__18328;
    wire N__18325;
    wire N__18322;
    wire N__18321;
    wire N__18320;
    wire N__18319;
    wire N__18318;
    wire N__18317;
    wire N__18314;
    wire N__18311;
    wire N__18308;
    wire N__18307;
    wire N__18306;
    wire N__18301;
    wire N__18294;
    wire N__18287;
    wire N__18280;
    wire N__18279;
    wire N__18278;
    wire N__18275;
    wire N__18274;
    wire N__18273;
    wire N__18272;
    wire N__18271;
    wire N__18270;
    wire N__18269;
    wire N__18264;
    wire N__18261;
    wire N__18254;
    wire N__18247;
    wire N__18238;
    wire N__18237;
    wire N__18236;
    wire N__18235;
    wire N__18234;
    wire N__18233;
    wire N__18232;
    wire N__18227;
    wire N__18226;
    wire N__18225;
    wire N__18224;
    wire N__18217;
    wire N__18212;
    wire N__18209;
    wire N__18204;
    wire N__18201;
    wire N__18190;
    wire N__18187;
    wire N__18186;
    wire N__18183;
    wire N__18180;
    wire N__18179;
    wire N__18176;
    wire N__18175;
    wire N__18174;
    wire N__18173;
    wire N__18172;
    wire N__18171;
    wire N__18168;
    wire N__18165;
    wire N__18162;
    wire N__18155;
    wire N__18152;
    wire N__18149;
    wire N__18146;
    wire N__18143;
    wire N__18130;
    wire N__18127;
    wire N__18124;
    wire N__18121;
    wire N__18118;
    wire N__18115;
    wire N__18112;
    wire N__18111;
    wire N__18108;
    wire N__18105;
    wire N__18102;
    wire N__18099;
    wire N__18096;
    wire N__18093;
    wire N__18088;
    wire N__18085;
    wire N__18084;
    wire N__18081;
    wire N__18078;
    wire N__18075;
    wire N__18070;
    wire N__18067;
    wire N__18064;
    wire N__18063;
    wire N__18062;
    wire N__18061;
    wire N__18060;
    wire N__18059;
    wire N__18058;
    wire N__18057;
    wire N__18056;
    wire N__18055;
    wire N__18054;
    wire N__18053;
    wire N__18048;
    wire N__18047;
    wire N__18046;
    wire N__18043;
    wire N__18042;
    wire N__18041;
    wire N__18038;
    wire N__18031;
    wire N__18026;
    wire N__18023;
    wire N__18018;
    wire N__18015;
    wire N__18014;
    wire N__18013;
    wire N__18010;
    wire N__18009;
    wire N__18008;
    wire N__18007;
    wire N__18006;
    wire N__18003;
    wire N__18000;
    wire N__17997;
    wire N__17994;
    wire N__17987;
    wire N__17982;
    wire N__17979;
    wire N__17976;
    wire N__17973;
    wire N__17966;
    wire N__17963;
    wire N__17960;
    wire N__17951;
    wire N__17946;
    wire N__17929;
    wire N__17928;
    wire N__17927;
    wire N__17926;
    wire N__17925;
    wire N__17924;
    wire N__17921;
    wire N__17920;
    wire N__17919;
    wire N__17918;
    wire N__17917;
    wire N__17916;
    wire N__17915;
    wire N__17914;
    wire N__17913;
    wire N__17912;
    wire N__17911;
    wire N__17910;
    wire N__17907;
    wire N__17906;
    wire N__17905;
    wire N__17904;
    wire N__17895;
    wire N__17894;
    wire N__17893;
    wire N__17892;
    wire N__17889;
    wire N__17888;
    wire N__17887;
    wire N__17886;
    wire N__17883;
    wire N__17876;
    wire N__17873;
    wire N__17870;
    wire N__17863;
    wire N__17862;
    wire N__17861;
    wire N__17860;
    wire N__17859;
    wire N__17856;
    wire N__17855;
    wire N__17854;
    wire N__17851;
    wire N__17848;
    wire N__17841;
    wire N__17838;
    wire N__17835;
    wire N__17832;
    wire N__17829;
    wire N__17828;
    wire N__17825;
    wire N__17818;
    wire N__17811;
    wire N__17806;
    wire N__17803;
    wire N__17800;
    wire N__17795;
    wire N__17792;
    wire N__17785;
    wire N__17778;
    wire N__17773;
    wire N__17770;
    wire N__17767;
    wire N__17760;
    wire N__17753;
    wire N__17750;
    wire N__17745;
    wire N__17742;
    wire N__17725;
    wire N__17724;
    wire N__17721;
    wire N__17718;
    wire N__17713;
    wire N__17710;
    wire N__17707;
    wire N__17704;
    wire N__17701;
    wire N__17698;
    wire N__17697;
    wire N__17696;
    wire N__17695;
    wire N__17694;
    wire N__17691;
    wire N__17688;
    wire N__17683;
    wire N__17680;
    wire N__17671;
    wire N__17668;
    wire N__17667;
    wire N__17664;
    wire N__17661;
    wire N__17660;
    wire N__17657;
    wire N__17654;
    wire N__17651;
    wire N__17650;
    wire N__17649;
    wire N__17642;
    wire N__17639;
    wire N__17636;
    wire N__17629;
    wire N__17626;
    wire N__17623;
    wire N__17620;
    wire N__17617;
    wire N__17616;
    wire N__17613;
    wire N__17610;
    wire N__17607;
    wire N__17602;
    wire N__17599;
    wire N__17596;
    wire N__17593;
    wire N__17590;
    wire N__17587;
    wire N__17584;
    wire N__17581;
    wire N__17578;
    wire N__17575;
    wire N__17572;
    wire N__17571;
    wire N__17568;
    wire N__17567;
    wire N__17566;
    wire N__17565;
    wire N__17562;
    wire N__17559;
    wire N__17554;
    wire N__17553;
    wire N__17552;
    wire N__17549;
    wire N__17548;
    wire N__17547;
    wire N__17546;
    wire N__17543;
    wire N__17538;
    wire N__17533;
    wire N__17532;
    wire N__17527;
    wire N__17526;
    wire N__17521;
    wire N__17516;
    wire N__17513;
    wire N__17510;
    wire N__17507;
    wire N__17504;
    wire N__17491;
    wire N__17488;
    wire N__17485;
    wire N__17482;
    wire N__17479;
    wire N__17476;
    wire N__17473;
    wire N__17472;
    wire N__17469;
    wire N__17466;
    wire N__17461;
    wire N__17458;
    wire N__17455;
    wire N__17452;
    wire N__17449;
    wire N__17446;
    wire N__17443;
    wire N__17442;
    wire N__17437;
    wire N__17434;
    wire N__17431;
    wire N__17428;
    wire N__17425;
    wire N__17422;
    wire N__17419;
    wire N__17416;
    wire N__17415;
    wire N__17412;
    wire N__17409;
    wire N__17404;
    wire N__17401;
    wire N__17398;
    wire N__17395;
    wire N__17394;
    wire N__17391;
    wire N__17388;
    wire N__17383;
    wire N__17380;
    wire N__17377;
    wire N__17374;
    wire N__17371;
    wire N__17368;
    wire N__17365;
    wire N__17364;
    wire N__17359;
    wire N__17356;
    wire N__17355;
    wire N__17352;
    wire N__17351;
    wire N__17350;
    wire N__17345;
    wire N__17340;
    wire N__17335;
    wire N__17332;
    wire N__17331;
    wire N__17328;
    wire N__17325;
    wire N__17322;
    wire N__17319;
    wire N__17316;
    wire N__17313;
    wire N__17308;
    wire N__17307;
    wire N__17306;
    wire N__17305;
    wire N__17304;
    wire N__17303;
    wire N__17302;
    wire N__17293;
    wire N__17290;
    wire N__17285;
    wire N__17282;
    wire N__17277;
    wire N__17274;
    wire N__17271;
    wire N__17266;
    wire N__17265;
    wire N__17264;
    wire N__17263;
    wire N__17262;
    wire N__17261;
    wire N__17260;
    wire N__17259;
    wire N__17258;
    wire N__17257;
    wire N__17254;
    wire N__17247;
    wire N__17244;
    wire N__17241;
    wire N__17232;
    wire N__17231;
    wire N__17230;
    wire N__17225;
    wire N__17222;
    wire N__17221;
    wire N__17216;
    wire N__17213;
    wire N__17210;
    wire N__17205;
    wire N__17202;
    wire N__17199;
    wire N__17194;
    wire N__17185;
    wire N__17184;
    wire N__17183;
    wire N__17182;
    wire N__17181;
    wire N__17178;
    wire N__17175;
    wire N__17172;
    wire N__17169;
    wire N__17166;
    wire N__17161;
    wire N__17156;
    wire N__17153;
    wire N__17148;
    wire N__17145;
    wire N__17142;
    wire N__17137;
    wire N__17134;
    wire N__17131;
    wire N__17128;
    wire N__17125;
    wire N__17122;
    wire N__17119;
    wire N__17116;
    wire N__17113;
    wire N__17112;
    wire N__17109;
    wire N__17106;
    wire N__17103;
    wire N__17100;
    wire N__17099;
    wire N__17094;
    wire N__17091;
    wire N__17088;
    wire N__17083;
    wire N__17080;
    wire N__17077;
    wire N__17074;
    wire N__17071;
    wire N__17068;
    wire N__17065;
    wire N__17062;
    wire N__17059;
    wire N__17056;
    wire N__17053;
    wire N__17050;
    wire N__17047;
    wire N__17044;
    wire N__17043;
    wire N__17042;
    wire N__17041;
    wire N__17040;
    wire N__17039;
    wire N__17038;
    wire N__17037;
    wire N__17034;
    wire N__17033;
    wire N__17032;
    wire N__17023;
    wire N__17012;
    wire N__17009;
    wire N__17002;
    wire N__17001;
    wire N__17000;
    wire N__16999;
    wire N__16998;
    wire N__16995;
    wire N__16994;
    wire N__16991;
    wire N__16988;
    wire N__16987;
    wire N__16984;
    wire N__16983;
    wire N__16980;
    wire N__16979;
    wire N__16970;
    wire N__16967;
    wire N__16958;
    wire N__16951;
    wire N__16948;
    wire N__16945;
    wire N__16942;
    wire N__16941;
    wire N__16940;
    wire N__16939;
    wire N__16938;
    wire N__16937;
    wire N__16936;
    wire N__16935;
    wire N__16934;
    wire N__16925;
    wire N__16922;
    wire N__16913;
    wire N__16906;
    wire N__16903;
    wire N__16900;
    wire N__16897;
    wire N__16894;
    wire N__16891;
    wire N__16888;
    wire N__16885;
    wire N__16882;
    wire N__16879;
    wire N__16876;
    wire N__16873;
    wire N__16870;
    wire N__16867;
    wire N__16864;
    wire N__16861;
    wire N__16858;
    wire N__16857;
    wire N__16852;
    wire N__16849;
    wire N__16846;
    wire N__16843;
    wire N__16840;
    wire N__16837;
    wire N__16834;
    wire N__16833;
    wire N__16828;
    wire N__16825;
    wire N__16822;
    wire N__16819;
    wire N__16816;
    wire N__16813;
    wire N__16810;
    wire N__16807;
    wire N__16804;
    wire N__16801;
    wire N__16798;
    wire N__16795;
    wire N__16792;
    wire N__16789;
    wire N__16788;
    wire N__16787;
    wire N__16786;
    wire N__16781;
    wire N__16780;
    wire N__16779;
    wire N__16778;
    wire N__16777;
    wire N__16772;
    wire N__16771;
    wire N__16770;
    wire N__16769;
    wire N__16768;
    wire N__16767;
    wire N__16764;
    wire N__16761;
    wire N__16758;
    wire N__16757;
    wire N__16756;
    wire N__16751;
    wire N__16748;
    wire N__16745;
    wire N__16740;
    wire N__16737;
    wire N__16734;
    wire N__16731;
    wire N__16728;
    wire N__16721;
    wire N__16702;
    wire N__16699;
    wire N__16696;
    wire N__16693;
    wire N__16690;
    wire N__16687;
    wire N__16684;
    wire N__16681;
    wire N__16678;
    wire N__16675;
    wire N__16672;
    wire N__16669;
    wire N__16666;
    wire N__16663;
    wire N__16660;
    wire N__16657;
    wire N__16654;
    wire N__16651;
    wire N__16648;
    wire N__16645;
    wire N__16644;
    wire N__16643;
    wire N__16642;
    wire N__16641;
    wire N__16640;
    wire N__16639;
    wire N__16636;
    wire N__16633;
    wire N__16628;
    wire N__16627;
    wire N__16622;
    wire N__16619;
    wire N__16618;
    wire N__16617;
    wire N__16616;
    wire N__16613;
    wire N__16608;
    wire N__16605;
    wire N__16604;
    wire N__16601;
    wire N__16598;
    wire N__16595;
    wire N__16590;
    wire N__16583;
    wire N__16580;
    wire N__16577;
    wire N__16564;
    wire N__16561;
    wire N__16558;
    wire N__16555;
    wire N__16552;
    wire N__16549;
    wire N__16546;
    wire N__16545;
    wire N__16544;
    wire N__16543;
    wire N__16540;
    wire N__16537;
    wire N__16534;
    wire N__16533;
    wire N__16530;
    wire N__16525;
    wire N__16520;
    wire N__16513;
    wire N__16512;
    wire N__16507;
    wire N__16506;
    wire N__16505;
    wire N__16504;
    wire N__16501;
    wire N__16500;
    wire N__16499;
    wire N__16498;
    wire N__16495;
    wire N__16492;
    wire N__16489;
    wire N__16486;
    wire N__16481;
    wire N__16478;
    wire N__16465;
    wire N__16462;
    wire N__16461;
    wire N__16458;
    wire N__16455;
    wire N__16452;
    wire N__16447;
    wire N__16446;
    wire N__16443;
    wire N__16442;
    wire N__16441;
    wire N__16440;
    wire N__16437;
    wire N__16434;
    wire N__16433;
    wire N__16430;
    wire N__16425;
    wire N__16422;
    wire N__16419;
    wire N__16416;
    wire N__16413;
    wire N__16402;
    wire N__16399;
    wire N__16398;
    wire N__16397;
    wire N__16392;
    wire N__16389;
    wire N__16388;
    wire N__16385;
    wire N__16380;
    wire N__16375;
    wire N__16374;
    wire N__16371;
    wire N__16368;
    wire N__16365;
    wire N__16364;
    wire N__16363;
    wire N__16362;
    wire N__16361;
    wire N__16358;
    wire N__16355;
    wire N__16346;
    wire N__16339;
    wire N__16336;
    wire N__16333;
    wire N__16332;
    wire N__16331;
    wire N__16330;
    wire N__16329;
    wire N__16326;
    wire N__16323;
    wire N__16316;
    wire N__16311;
    wire N__16306;
    wire N__16303;
    wire N__16300;
    wire N__16297;
    wire N__16294;
    wire N__16291;
    wire N__16288;
    wire N__16285;
    wire N__16282;
    wire N__16279;
    wire N__16276;
    wire N__16275;
    wire N__16274;
    wire N__16273;
    wire N__16272;
    wire N__16271;
    wire N__16268;
    wire N__16267;
    wire N__16260;
    wire N__16259;
    wire N__16258;
    wire N__16257;
    wire N__16256;
    wire N__16255;
    wire N__16254;
    wire N__16253;
    wire N__16252;
    wire N__16251;
    wire N__16250;
    wire N__16247;
    wire N__16244;
    wire N__16241;
    wire N__16238;
    wire N__16235;
    wire N__16232;
    wire N__16227;
    wire N__16218;
    wire N__16209;
    wire N__16192;
    wire N__16189;
    wire N__16186;
    wire N__16183;
    wire N__16180;
    wire N__16177;
    wire N__16174;
    wire N__16173;
    wire N__16172;
    wire N__16169;
    wire N__16164;
    wire N__16159;
    wire N__16156;
    wire N__16155;
    wire N__16152;
    wire N__16151;
    wire N__16150;
    wire N__16147;
    wire N__16144;
    wire N__16137;
    wire N__16132;
    wire N__16131;
    wire N__16130;
    wire N__16129;
    wire N__16122;
    wire N__16121;
    wire N__16120;
    wire N__16119;
    wire N__16118;
    wire N__16115;
    wire N__16112;
    wire N__16111;
    wire N__16110;
    wire N__16109;
    wire N__16108;
    wire N__16105;
    wire N__16104;
    wire N__16103;
    wire N__16098;
    wire N__16095;
    wire N__16092;
    wire N__16089;
    wire N__16084;
    wire N__16081;
    wire N__16072;
    wire N__16057;
    wire N__16054;
    wire N__16053;
    wire N__16052;
    wire N__16047;
    wire N__16044;
    wire N__16041;
    wire N__16038;
    wire N__16033;
    wire N__16030;
    wire N__16029;
    wire N__16026;
    wire N__16023;
    wire N__16020;
    wire N__16015;
    wire N__16012;
    wire N__16009;
    wire N__16006;
    wire N__16005;
    wire N__16004;
    wire N__16001;
    wire N__15996;
    wire N__15993;
    wire N__15988;
    wire N__15985;
    wire N__15982;
    wire N__15979;
    wire N__15978;
    wire N__15977;
    wire N__15976;
    wire N__15975;
    wire N__15974;
    wire N__15973;
    wire N__15972;
    wire N__15955;
    wire N__15954;
    wire N__15951;
    wire N__15948;
    wire N__15943;
    wire N__15942;
    wire N__15941;
    wire N__15938;
    wire N__15935;
    wire N__15932;
    wire N__15931;
    wire N__15930;
    wire N__15929;
    wire N__15928;
    wire N__15927;
    wire N__15926;
    wire N__15925;
    wire N__15924;
    wire N__15923;
    wire N__15922;
    wire N__15921;
    wire N__15920;
    wire N__15919;
    wire N__15902;
    wire N__15897;
    wire N__15892;
    wire N__15887;
    wire N__15882;
    wire N__15871;
    wire N__15870;
    wire N__15867;
    wire N__15864;
    wire N__15861;
    wire N__15858;
    wire N__15855;
    wire N__15852;
    wire N__15849;
    wire N__15844;
    wire N__15843;
    wire N__15842;
    wire N__15839;
    wire N__15838;
    wire N__15837;
    wire N__15836;
    wire N__15835;
    wire N__15832;
    wire N__15829;
    wire N__15826;
    wire N__15817;
    wire N__15814;
    wire N__15805;
    wire N__15804;
    wire N__15803;
    wire N__15800;
    wire N__15797;
    wire N__15796;
    wire N__15795;
    wire N__15794;
    wire N__15793;
    wire N__15790;
    wire N__15787;
    wire N__15784;
    wire N__15781;
    wire N__15778;
    wire N__15773;
    wire N__15760;
    wire N__15757;
    wire N__15754;
    wire N__15751;
    wire N__15748;
    wire N__15745;
    wire N__15744;
    wire N__15741;
    wire N__15740;
    wire N__15737;
    wire N__15730;
    wire N__15727;
    wire N__15724;
    wire N__15721;
    wire N__15720;
    wire N__15717;
    wire N__15712;
    wire N__15709;
    wire N__15706;
    wire N__15703;
    wire N__15700;
    wire N__15699;
    wire N__15696;
    wire N__15691;
    wire N__15688;
    wire N__15685;
    wire N__15682;
    wire N__15681;
    wire N__15676;
    wire N__15673;
    wire N__15670;
    wire N__15669;
    wire N__15666;
    wire N__15663;
    wire N__15658;
    wire N__15655;
    wire N__15652;
    wire N__15649;
    wire N__15646;
    wire N__15643;
    wire N__15640;
    wire N__15637;
    wire N__15636;
    wire N__15633;
    wire N__15630;
    wire N__15625;
    wire N__15624;
    wire N__15621;
    wire N__15620;
    wire N__15619;
    wire N__15616;
    wire N__15613;
    wire N__15608;
    wire N__15601;
    wire N__15598;
    wire N__15595;
    wire N__15592;
    wire N__15589;
    wire N__15586;
    wire N__15583;
    wire N__15582;
    wire N__15579;
    wire N__15576;
    wire N__15575;
    wire N__15572;
    wire N__15569;
    wire N__15568;
    wire N__15565;
    wire N__15562;
    wire N__15559;
    wire N__15554;
    wire N__15551;
    wire N__15544;
    wire N__15541;
    wire N__15538;
    wire N__15537;
    wire N__15534;
    wire N__15531;
    wire N__15528;
    wire N__15525;
    wire N__15522;
    wire N__15517;
    wire N__15514;
    wire N__15513;
    wire N__15510;
    wire N__15507;
    wire N__15504;
    wire N__15501;
    wire N__15496;
    wire N__15493;
    wire N__15490;
    wire N__15487;
    wire N__15484;
    wire N__15483;
    wire N__15482;
    wire N__15481;
    wire N__15480;
    wire N__15477;
    wire N__15476;
    wire N__15475;
    wire N__15474;
    wire N__15473;
    wire N__15472;
    wire N__15467;
    wire N__15462;
    wire N__15459;
    wire N__15456;
    wire N__15451;
    wire N__15446;
    wire N__15443;
    wire N__15440;
    wire N__15435;
    wire N__15434;
    wire N__15429;
    wire N__15424;
    wire N__15421;
    wire N__15418;
    wire N__15409;
    wire N__15406;
    wire N__15403;
    wire N__15400;
    wire N__15397;
    wire N__15394;
    wire N__15391;
    wire N__15388;
    wire N__15385;
    wire N__15384;
    wire N__15381;
    wire N__15378;
    wire N__15377;
    wire N__15374;
    wire N__15371;
    wire N__15368;
    wire N__15363;
    wire N__15358;
    wire N__15357;
    wire N__15352;
    wire N__15349;
    wire N__15346;
    wire N__15343;
    wire N__15340;
    wire N__15337;
    wire N__15336;
    wire N__15333;
    wire N__15330;
    wire N__15327;
    wire N__15324;
    wire N__15321;
    wire N__15320;
    wire N__15317;
    wire N__15314;
    wire N__15311;
    wire N__15304;
    wire N__15301;
    wire N__15298;
    wire N__15297;
    wire N__15294;
    wire N__15291;
    wire N__15286;
    wire N__15283;
    wire N__15280;
    wire N__15279;
    wire N__15276;
    wire N__15273;
    wire N__15268;
    wire N__15265;
    wire N__15262;
    wire N__15259;
    wire N__15256;
    wire N__15253;
    wire N__15250;
    wire N__15247;
    wire N__15244;
    wire N__15241;
    wire N__15238;
    wire N__15235;
    wire N__15232;
    wire N__15229;
    wire N__15226;
    wire N__15223;
    wire N__15220;
    wire N__15217;
    wire N__15214;
    wire N__15211;
    wire N__15208;
    wire N__15205;
    wire N__15202;
    wire N__15199;
    wire N__15196;
    wire N__15193;
    wire N__15192;
    wire N__15189;
    wire N__15186;
    wire N__15181;
    wire N__15178;
    wire N__15175;
    wire N__15172;
    wire N__15169;
    wire N__15166;
    wire N__15163;
    wire N__15160;
    wire N__15157;
    wire N__15154;
    wire N__15151;
    wire N__15148;
    wire N__15145;
    wire N__15142;
    wire N__15139;
    wire N__15136;
    wire N__15133;
    wire N__15130;
    wire N__15127;
    wire N__15126;
    wire N__15121;
    wire N__15118;
    wire N__15117;
    wire N__15112;
    wire N__15111;
    wire N__15110;
    wire N__15109;
    wire N__15108;
    wire N__15107;
    wire N__15104;
    wire N__15099;
    wire N__15096;
    wire N__15091;
    wire N__15088;
    wire N__15081;
    wire N__15076;
    wire N__15073;
    wire N__15072;
    wire N__15067;
    wire N__15064;
    wire N__15061;
    wire N__15060;
    wire N__15059;
    wire N__15056;
    wire N__15055;
    wire N__15050;
    wire N__15047;
    wire N__15044;
    wire N__15041;
    wire N__15040;
    wire N__15039;
    wire N__15038;
    wire N__15035;
    wire N__15032;
    wire N__15029;
    wire N__15022;
    wire N__15013;
    wire N__15010;
    wire N__15007;
    wire N__15004;
    wire N__15001;
    wire N__15000;
    wire N__14995;
    wire N__14992;
    wire N__14989;
    wire N__14986;
    wire N__14983;
    wire N__14980;
    wire N__14977;
    wire N__14974;
    wire N__14971;
    wire N__14968;
    wire N__14965;
    wire N__14962;
    wire N__14959;
    wire N__14956;
    wire N__14953;
    wire N__14950;
    wire N__14947;
    wire N__14944;
    wire N__14941;
    wire N__14938;
    wire N__14935;
    wire N__14932;
    wire N__14929;
    wire N__14926;
    wire N__14923;
    wire N__14920;
    wire N__14919;
    wire N__14918;
    wire N__14917;
    wire N__14910;
    wire N__14909;
    wire N__14908;
    wire N__14907;
    wire N__14906;
    wire N__14903;
    wire N__14900;
    wire N__14899;
    wire N__14898;
    wire N__14891;
    wire N__14888;
    wire N__14885;
    wire N__14882;
    wire N__14877;
    wire N__14874;
    wire N__14863;
    wire N__14860;
    wire N__14857;
    wire N__14854;
    wire N__14851;
    wire N__14848;
    wire N__14845;
    wire N__14842;
    wire N__14841;
    wire N__14840;
    wire N__14839;
    wire N__14838;
    wire N__14837;
    wire N__14836;
    wire N__14835;
    wire N__14826;
    wire N__14817;
    wire N__14812;
    wire N__14811;
    wire N__14810;
    wire N__14809;
    wire N__14808;
    wire N__14805;
    wire N__14804;
    wire N__14803;
    wire N__14800;
    wire N__14797;
    wire N__14796;
    wire N__14795;
    wire N__14786;
    wire N__14777;
    wire N__14774;
    wire N__14767;
    wire N__14766;
    wire N__14765;
    wire N__14764;
    wire N__14763;
    wire N__14762;
    wire N__14761;
    wire N__14758;
    wire N__14755;
    wire N__14754;
    wire N__14751;
    wire N__14742;
    wire N__14733;
    wire N__14728;
    wire N__14727;
    wire N__14724;
    wire N__14721;
    wire N__14720;
    wire N__14719;
    wire N__14718;
    wire N__14717;
    wire N__14716;
    wire N__14715;
    wire N__14706;
    wire N__14697;
    wire N__14692;
    wire N__14689;
    wire N__14686;
    wire N__14683;
    wire N__14680;
    wire N__14677;
    wire N__14674;
    wire N__14671;
    wire N__14668;
    wire N__14665;
    wire N__14662;
    wire N__14659;
    wire N__14656;
    wire N__14653;
    wire N__14650;
    wire N__14647;
    wire N__14644;
    wire N__14641;
    wire N__14640;
    wire N__14635;
    wire N__14632;
    wire N__14629;
    wire N__14626;
    wire N__14623;
    wire N__14620;
    wire N__14617;
    wire N__14614;
    wire N__14611;
    wire N__14608;
    wire N__14605;
    wire N__14602;
    wire N__14599;
    wire N__14596;
    wire N__14593;
    wire N__14590;
    wire N__14589;
    wire N__14586;
    wire N__14585;
    wire N__14578;
    wire N__14575;
    wire N__14572;
    wire N__14569;
    wire N__14566;
    wire N__14563;
    wire N__14560;
    wire N__14557;
    wire N__14554;
    wire N__14551;
    wire N__14548;
    wire N__14545;
    wire N__14542;
    wire N__14539;
    wire N__14536;
    wire N__14533;
    wire N__14530;
    wire N__14527;
    wire N__14524;
    wire N__14521;
    wire N__14518;
    wire N__14515;
    wire N__14512;
    wire N__14509;
    wire N__14508;
    wire N__14505;
    wire N__14502;
    wire N__14501;
    wire N__14500;
    wire N__14497;
    wire N__14494;
    wire N__14491;
    wire N__14488;
    wire N__14483;
    wire N__14480;
    wire N__14477;
    wire N__14474;
    wire N__14467;
    wire N__14464;
    wire N__14461;
    wire N__14458;
    wire N__14455;
    wire N__14452;
    wire N__14449;
    wire N__14446;
    wire N__14443;
    wire N__14440;
    wire N__14437;
    wire N__14434;
    wire N__14431;
    wire N__14428;
    wire N__14427;
    wire N__14424;
    wire N__14421;
    wire N__14416;
    wire N__14415;
    wire N__14414;
    wire N__14413;
    wire N__14410;
    wire N__14407;
    wire N__14402;
    wire N__14395;
    wire N__14392;
    wire N__14389;
    wire N__14386;
    wire N__14383;
    wire N__14380;
    wire N__14379;
    wire N__14376;
    wire N__14375;
    wire N__14372;
    wire N__14367;
    wire N__14362;
    wire N__14361;
    wire N__14358;
    wire N__14353;
    wire N__14350;
    wire N__14347;
    wire N__14344;
    wire N__14341;
    wire N__14338;
    wire N__14335;
    wire N__14332;
    wire N__14329;
    wire N__14328;
    wire N__14323;
    wire N__14320;
    wire N__14317;
    wire N__14314;
    wire N__14313;
    wire N__14308;
    wire N__14305;
    wire N__14304;
    wire N__14299;
    wire N__14296;
    wire N__14293;
    wire N__14292;
    wire N__14289;
    wire N__14286;
    wire N__14283;
    wire N__14278;
    wire N__14275;
    wire N__14272;
    wire N__14269;
    wire N__14268;
    wire N__14265;
    wire N__14262;
    wire N__14259;
    wire N__14256;
    wire N__14253;
    wire N__14250;
    wire N__14247;
    wire N__14242;
    wire N__14239;
    wire N__14236;
    wire N__14233;
    wire N__14230;
    wire N__14227;
    wire N__14224;
    wire N__14223;
    wire N__14222;
    wire N__14219;
    wire N__14214;
    wire N__14209;
    wire N__14206;
    wire N__14205;
    wire N__14202;
    wire N__14199;
    wire N__14194;
    wire N__14191;
    wire N__14188;
    wire N__14185;
    wire N__14182;
    wire N__14179;
    wire N__14176;
    wire N__14175;
    wire N__14172;
    wire N__14169;
    wire N__14164;
    wire N__14161;
    wire N__14160;
    wire N__14157;
    wire N__14156;
    wire N__14153;
    wire N__14150;
    wire N__14147;
    wire N__14140;
    wire N__14137;
    wire N__14134;
    wire N__14131;
    wire N__14128;
    wire N__14125;
    wire N__14122;
    wire N__14119;
    wire N__14116;
    wire N__14113;
    wire N__14110;
    wire N__14107;
    wire N__14104;
    wire N__14101;
    wire N__14098;
    wire N__14097;
    wire N__14096;
    wire N__14095;
    wire N__14092;
    wire N__14089;
    wire N__14088;
    wire N__14087;
    wire N__14084;
    wire N__14083;
    wire N__14080;
    wire N__14077;
    wire N__14064;
    wire N__14059;
    wire N__14056;
    wire N__14053;
    wire N__14050;
    wire N__14047;
    wire N__14044;
    wire N__14041;
    wire N__14038;
    wire N__14035;
    wire N__14034;
    wire N__14033;
    wire N__14026;
    wire N__14025;
    wire N__14022;
    wire N__14019;
    wire N__14016;
    wire N__14011;
    wire N__14008;
    wire N__14007;
    wire N__14004;
    wire N__14001;
    wire N__13998;
    wire N__13995;
    wire N__13992;
    wire N__13987;
    wire N__13984;
    wire N__13981;
    wire N__13978;
    wire N__13975;
    wire N__13974;
    wire N__13971;
    wire N__13968;
    wire N__13965;
    wire N__13962;
    wire N__13957;
    wire N__13954;
    wire N__13951;
    wire N__13948;
    wire N__13945;
    wire N__13942;
    wire N__13939;
    wire N__13938;
    wire N__13935;
    wire N__13932;
    wire N__13929;
    wire N__13926;
    wire N__13921;
    wire N__13920;
    wire N__13917;
    wire N__13914;
    wire N__13909;
    wire N__13906;
    wire N__13903;
    wire N__13900;
    wire N__13897;
    wire N__13896;
    wire N__13893;
    wire N__13890;
    wire N__13887;
    wire N__13884;
    wire N__13881;
    wire N__13878;
    wire N__13873;
    wire N__13870;
    wire N__13867;
    wire N__13864;
    wire N__13863;
    wire N__13862;
    wire N__13859;
    wire N__13854;
    wire N__13851;
    wire N__13848;
    wire N__13845;
    wire N__13842;
    wire N__13837;
    wire N__13834;
    wire N__13831;
    wire N__13830;
    wire N__13829;
    wire N__13824;
    wire N__13821;
    wire N__13818;
    wire N__13815;
    wire N__13812;
    wire N__13809;
    wire N__13804;
    wire N__13801;
    wire N__13798;
    wire N__13795;
    wire N__13792;
    wire N__13789;
    wire N__13786;
    wire N__13783;
    wire N__13780;
    wire N__13777;
    wire N__13774;
    wire N__13771;
    wire N__13768;
    wire N__13765;
    wire N__13762;
    wire N__13759;
    wire N__13756;
    wire N__13753;
    wire N__13750;
    wire N__13747;
    wire N__13744;
    wire N__13741;
    wire N__13738;
    wire N__13735;
    wire N__13732;
    wire N__13729;
    wire N__13726;
    wire N__13725;
    wire N__13722;
    wire N__13719;
    wire N__13714;
    wire N__13711;
    wire N__13708;
    wire N__13705;
    wire N__13702;
    wire N__13699;
    wire N__13696;
    wire N__13693;
    wire N__13692;
    wire N__13689;
    wire N__13688;
    wire N__13685;
    wire N__13684;
    wire N__13681;
    wire N__13674;
    wire N__13669;
    wire N__13666;
    wire N__13663;
    wire N__13662;
    wire N__13659;
    wire N__13656;
    wire N__13655;
    wire N__13654;
    wire N__13651;
    wire N__13648;
    wire N__13643;
    wire N__13636;
    wire N__13633;
    wire N__13630;
    wire N__13627;
    wire N__13626;
    wire N__13625;
    wire N__13624;
    wire N__13623;
    wire N__13620;
    wire N__13615;
    wire N__13610;
    wire N__13603;
    wire N__13600;
    wire N__13597;
    wire N__13594;
    wire N__13593;
    wire N__13590;
    wire N__13589;
    wire N__13586;
    wire N__13585;
    wire N__13584;
    wire N__13583;
    wire N__13580;
    wire N__13573;
    wire N__13568;
    wire N__13561;
    wire N__13558;
    wire N__13557;
    wire N__13556;
    wire N__13553;
    wire N__13550;
    wire N__13547;
    wire N__13544;
    wire N__13539;
    wire N__13534;
    wire N__13531;
    wire N__13528;
    wire N__13525;
    wire N__13522;
    wire N__13519;
    wire N__13516;
    wire N__13513;
    wire N__13510;
    wire N__13507;
    wire N__13504;
    wire N__13501;
    wire N__13498;
    wire N__13495;
    wire N__13492;
    wire N__13489;
    wire N__13486;
    wire N__13483;
    wire N__13480;
    wire N__13477;
    wire N__13474;
    wire N__13471;
    wire N__13468;
    wire N__13467;
    wire N__13466;
    wire N__13463;
    wire N__13460;
    wire N__13457;
    wire N__13454;
    wire N__13451;
    wire N__13450;
    wire N__13447;
    wire N__13444;
    wire N__13441;
    wire N__13438;
    wire N__13435;
    wire N__13426;
    wire N__13425;
    wire N__13422;
    wire N__13419;
    wire N__13416;
    wire N__13411;
    wire N__13408;
    wire N__13407;
    wire N__13402;
    wire N__13399;
    wire N__13396;
    wire N__13393;
    wire N__13390;
    wire N__13387;
    wire N__13384;
    wire N__13383;
    wire N__13380;
    wire N__13377;
    wire N__13372;
    wire N__13369;
    wire N__13366;
    wire N__13363;
    wire N__13360;
    wire N__13357;
    wire N__13356;
    wire N__13355;
    wire N__13352;
    wire N__13349;
    wire N__13346;
    wire N__13339;
    wire N__13336;
    wire N__13333;
    wire N__13330;
    wire N__13329;
    wire N__13326;
    wire N__13321;
    wire N__13318;
    wire N__13315;
    wire N__13312;
    wire N__13309;
    wire N__13308;
    wire N__13307;
    wire N__13300;
    wire N__13297;
    wire N__13296;
    wire N__13293;
    wire N__13292;
    wire N__13285;
    wire N__13282;
    wire N__13279;
    wire N__13276;
    wire N__13273;
    wire N__13270;
    wire N__13267;
    wire N__13264;
    wire N__13261;
    wire N__13258;
    wire N__13255;
    wire N__13252;
    wire N__13249;
    wire N__13246;
    wire N__13243;
    wire N__13240;
    wire N__13237;
    wire N__13234;
    wire N__13233;
    wire N__13230;
    wire N__13227;
    wire N__13224;
    wire N__13223;
    wire N__13220;
    wire N__13217;
    wire N__13216;
    wire N__13213;
    wire N__13210;
    wire N__13207;
    wire N__13204;
    wire N__13195;
    wire N__13192;
    wire N__13191;
    wire N__13186;
    wire N__13183;
    wire N__13182;
    wire N__13177;
    wire N__13174;
    wire N__13171;
    wire N__13168;
    wire N__13167;
    wire N__13162;
    wire N__13159;
    wire N__13156;
    wire N__13153;
    wire N__13150;
    wire N__13147;
    wire N__13144;
    wire N__13141;
    wire N__13138;
    wire N__13135;
    wire N__13132;
    wire N__13129;
    wire N__13126;
    wire N__13123;
    wire N__13120;
    wire N__13117;
    wire N__13116;
    wire N__13115;
    wire N__13114;
    wire N__13113;
    wire N__13106;
    wire N__13103;
    wire N__13100;
    wire N__13097;
    wire N__13090;
    wire N__13089;
    wire N__13088;
    wire N__13085;
    wire N__13080;
    wire N__13079;
    wire N__13078;
    wire N__13077;
    wire N__13074;
    wire N__13071;
    wire N__13066;
    wire N__13063;
    wire N__13060;
    wire N__13057;
    wire N__13048;
    wire N__13045;
    wire N__13044;
    wire N__13039;
    wire N__13036;
    wire N__13033;
    wire N__13030;
    wire N__13027;
    wire N__13024;
    wire N__13023;
    wire N__13018;
    wire N__13015;
    wire N__13012;
    wire N__13011;
    wire N__13008;
    wire N__13007;
    wire N__13004;
    wire N__13001;
    wire N__12998;
    wire N__12995;
    wire N__12990;
    wire N__12989;
    wire N__12988;
    wire N__12987;
    wire N__12986;
    wire N__12985;
    wire N__12984;
    wire N__12983;
    wire N__12982;
    wire N__12981;
    wire N__12978;
    wire N__12975;
    wire N__12968;
    wire N__12963;
    wire N__12954;
    wire N__12951;
    wire N__12940;
    wire N__12939;
    wire N__12938;
    wire N__12935;
    wire N__12932;
    wire N__12929;
    wire N__12926;
    wire N__12919;
    wire N__12916;
    wire N__12915;
    wire N__12912;
    wire N__12909;
    wire N__12906;
    wire N__12903;
    wire N__12900;
    wire N__12897;
    wire N__12892;
    wire N__12889;
    wire N__12886;
    wire N__12883;
    wire N__12880;
    wire N__12877;
    wire N__12874;
    wire N__12871;
    wire N__12870;
    wire N__12865;
    wire N__12862;
    wire N__12859;
    wire N__12856;
    wire N__12853;
    wire N__12850;
    wire N__12847;
    wire N__12844;
    wire N__12841;
    wire N__12838;
    wire N__12835;
    wire N__12832;
    wire N__12831;
    wire N__12830;
    wire N__12827;
    wire N__12826;
    wire N__12825;
    wire N__12820;
    wire N__12819;
    wire N__12818;
    wire N__12817;
    wire N__12816;
    wire N__12815;
    wire N__12814;
    wire N__12813;
    wire N__12812;
    wire N__12811;
    wire N__12808;
    wire N__12803;
    wire N__12800;
    wire N__12799;
    wire N__12798;
    wire N__12781;
    wire N__12778;
    wire N__12771;
    wire N__12766;
    wire N__12757;
    wire N__12754;
    wire N__12751;
    wire N__12748;
    wire N__12745;
    wire N__12742;
    wire N__12739;
    wire N__12736;
    wire N__12733;
    wire N__12730;
    wire N__12729;
    wire N__12726;
    wire N__12723;
    wire N__12720;
    wire N__12717;
    wire N__12712;
    wire N__12709;
    wire N__12706;
    wire N__12703;
    wire N__12700;
    wire N__12697;
    wire N__12694;
    wire N__12691;
    wire N__12688;
    wire N__12685;
    wire N__12682;
    wire N__12679;
    wire N__12676;
    wire N__12673;
    wire N__12670;
    wire N__12667;
    wire N__12666;
    wire N__12661;
    wire N__12658;
    wire N__12655;
    wire N__12652;
    wire N__12649;
    wire N__12646;
    wire N__12643;
    wire N__12640;
    wire N__12637;
    wire N__12634;
    wire N__12631;
    wire N__12628;
    wire N__12625;
    wire N__12622;
    wire N__12619;
    wire N__12616;
    wire N__12613;
    wire N__12610;
    wire N__12609;
    wire N__12606;
    wire N__12603;
    wire N__12600;
    wire N__12595;
    wire N__12592;
    wire N__12589;
    wire N__12586;
    wire N__12583;
    wire N__12580;
    wire N__12577;
    wire N__12574;
    wire N__12571;
    wire N__12568;
    wire N__12565;
    wire N__12562;
    wire N__12559;
    wire N__12556;
    wire N__12553;
    wire N__12550;
    wire N__12547;
    wire N__12544;
    wire N__12541;
    wire N__12538;
    wire N__12535;
    wire N__12532;
    wire N__12529;
    wire N__12526;
    wire N__12525;
    wire N__12524;
    wire N__12523;
    wire N__12514;
    wire N__12513;
    wire N__12512;
    wire N__12509;
    wire N__12506;
    wire N__12503;
    wire N__12498;
    wire N__12493;
    wire N__12490;
    wire N__12487;
    wire N__12484;
    wire N__12481;
    wire N__12480;
    wire N__12475;
    wire N__12474;
    wire N__12473;
    wire N__12470;
    wire N__12467;
    wire N__12464;
    wire N__12461;
    wire N__12458;
    wire N__12451;
    wire N__12450;
    wire N__12449;
    wire N__12446;
    wire N__12441;
    wire N__12438;
    wire N__12433;
    wire N__12430;
    wire N__12427;
    wire N__12426;
    wire N__12423;
    wire N__12420;
    wire N__12417;
    wire N__12412;
    wire N__12411;
    wire N__12406;
    wire N__12403;
    wire N__12402;
    wire N__12401;
    wire N__12400;
    wire N__12397;
    wire N__12394;
    wire N__12389;
    wire N__12382;
    wire N__12379;
    wire N__12376;
    wire N__12375;
    wire N__12374;
    wire N__12373;
    wire N__12370;
    wire N__12367;
    wire N__12364;
    wire N__12361;
    wire N__12358;
    wire N__12355;
    wire N__12346;
    wire N__12345;
    wire N__12344;
    wire N__12343;
    wire N__12342;
    wire N__12331;
    wire N__12328;
    wire N__12325;
    wire N__12322;
    wire N__12319;
    wire N__12316;
    wire N__12313;
    wire N__12310;
    wire N__12307;
    wire N__12304;
    wire N__12301;
    wire N__12298;
    wire N__12295;
    wire N__12292;
    wire N__12289;
    wire N__12286;
    wire N__12283;
    wire N__12280;
    wire N__12277;
    wire N__12274;
    wire N__12271;
    wire N__12268;
    wire N__12265;
    wire N__12262;
    wire N__12259;
    wire N__12256;
    wire N__12253;
    wire N__12250;
    wire N__12247;
    wire N__12244;
    wire N__12241;
    wire N__12238;
    wire N__12235;
    wire N__12232;
    wire N__12229;
    wire N__12226;
    wire N__12223;
    wire N__12220;
    wire N__12217;
    wire N__12214;
    wire N__12211;
    wire N__12208;
    wire N__12205;
    wire N__12202;
    wire N__12201;
    wire N__12200;
    wire N__12199;
    wire N__12198;
    wire N__12187;
    wire N__12184;
    wire N__12183;
    wire N__12182;
    wire N__12181;
    wire N__12178;
    wire N__12177;
    wire N__12172;
    wire N__12165;
    wire N__12160;
    wire N__12159;
    wire N__12158;
    wire N__12155;
    wire N__12148;
    wire N__12145;
    wire N__12142;
    wire N__12139;
    wire N__12136;
    wire N__12133;
    wire N__12130;
    wire N__12127;
    wire N__12126;
    wire N__12125;
    wire N__12124;
    wire N__12123;
    wire N__12112;
    wire N__12109;
    wire N__12108;
    wire N__12107;
    wire N__12100;
    wire N__12097;
    wire N__12094;
    wire N__12091;
    wire N__12088;
    wire N__12085;
    wire N__12082;
    wire N__12079;
    wire N__12078;
    wire N__12077;
    wire N__12074;
    wire N__12071;
    wire N__12068;
    wire N__12065;
    wire N__12058;
    wire N__12057;
    wire N__12056;
    wire N__12053;
    wire N__12048;
    wire N__12043;
    wire N__12042;
    wire N__12039;
    wire N__12036;
    wire N__12031;
    wire N__12028;
    wire N__12025;
    wire N__12024;
    wire N__12023;
    wire N__12022;
    wire N__12019;
    wire N__12012;
    wire N__12007;
    wire N__12006;
    wire N__12005;
    wire N__12000;
    wire N__11997;
    wire N__11992;
    wire N__11989;
    wire N__11986;
    wire N__11983;
    wire N__11980;
    wire N__11977;
    wire N__11974;
    wire N__11971;
    wire N__11968;
    wire N__11965;
    wire N__11962;
    wire N__11959;
    wire N__11956;
    wire N__11953;
    wire N__11950;
    wire N__11947;
    wire N__11944;
    wire N__11941;
    wire N__11938;
    wire N__11935;
    wire N__11932;
    wire N__11929;
    wire N__11926;
    wire N__11923;
    wire N__11920;
    wire N__11917;
    wire N__11914;
    wire N__11911;
    wire N__11908;
    wire N__11905;
    wire N__11902;
    wire N__11899;
    wire N__11896;
    wire N__11893;
    wire N__11890;
    wire N__11887;
    wire N__11884;
    wire N__11881;
    wire N__11878;
    wire N__11875;
    wire N__11872;
    wire N__11871;
    wire N__11870;
    wire N__11869;
    wire N__11868;
    wire N__11857;
    wire N__11854;
    wire N__11853;
    wire N__11852;
    wire N__11849;
    wire N__11846;
    wire N__11839;
    wire N__11836;
    wire N__11835;
    wire N__11834;
    wire N__11831;
    wire N__11830;
    wire N__11823;
    wire N__11820;
    wire N__11815;
    wire N__11814;
    wire N__11811;
    wire N__11808;
    wire N__11803;
    wire N__11802;
    wire N__11801;
    wire N__11798;
    wire N__11793;
    wire N__11790;
    wire N__11785;
    wire N__11782;
    wire N__11779;
    wire N__11776;
    wire N__11773;
    wire N__11770;
    wire N__11767;
    wire N__11764;
    wire N__11761;
    wire N__11758;
    wire N__11755;
    wire N__11752;
    wire N__11749;
    wire N__11746;
    wire N__11743;
    wire N__11740;
    wire N__11737;
    wire N__11736;
    wire N__11735;
    wire N__11734;
    wire N__11733;
    wire N__11732;
    wire N__11729;
    wire N__11726;
    wire N__11725;
    wire N__11724;
    wire N__11723;
    wire N__11720;
    wire N__11717;
    wire N__11716;
    wire N__11709;
    wire N__11706;
    wire N__11699;
    wire N__11692;
    wire N__11683;
    wire N__11682;
    wire N__11681;
    wire N__11676;
    wire N__11673;
    wire N__11670;
    wire N__11665;
    wire N__11662;
    wire N__11661;
    wire N__11660;
    wire N__11659;
    wire N__11654;
    wire N__11649;
    wire N__11644;
    wire N__11641;
    wire N__11640;
    wire N__11639;
    wire N__11638;
    wire N__11637;
    wire N__11630;
    wire N__11625;
    wire N__11620;
    wire N__11617;
    wire N__11616;
    wire N__11615;
    wire N__11608;
    wire N__11605;
    wire N__11604;
    wire N__11603;
    wire N__11600;
    wire N__11593;
    wire N__11590;
    wire N__11589;
    wire N__11588;
    wire N__11583;
    wire N__11580;
    wire N__11575;
    wire N__11572;
    wire N__11569;
    wire N__11566;
    wire N__11565;
    wire N__11564;
    wire N__11563;
    wire N__11560;
    wire N__11557;
    wire N__11554;
    wire N__11551;
    wire N__11550;
    wire N__11547;
    wire N__11544;
    wire N__11537;
    wire N__11530;
    wire N__11527;
    wire N__11526;
    wire N__11525;
    wire N__11524;
    wire N__11523;
    wire N__11520;
    wire N__11519;
    wire N__11518;
    wire N__11517;
    wire N__11516;
    wire N__11513;
    wire N__11506;
    wire N__11503;
    wire N__11494;
    wire N__11491;
    wire N__11482;
    wire N__11481;
    wire N__11480;
    wire N__11477;
    wire N__11474;
    wire N__11471;
    wire N__11468;
    wire N__11465;
    wire N__11458;
    wire N__11457;
    wire N__11456;
    wire N__11455;
    wire N__11452;
    wire N__11445;
    wire N__11442;
    wire N__11437;
    wire N__11434;
    wire N__11431;
    wire N__11428;
    wire N__11425;
    wire N__11422;
    wire N__11419;
    wire N__11418;
    wire N__11415;
    wire N__11414;
    wire N__11409;
    wire N__11406;
    wire N__11401;
    wire N__11398;
    wire N__11397;
    wire N__11396;
    wire N__11395;
    wire N__11386;
    wire N__11383;
    wire N__11382;
    wire N__11381;
    wire N__11380;
    wire N__11375;
    wire N__11370;
    wire N__11365;
    wire N__11362;
    wire N__11361;
    wire N__11360;
    wire N__11357;
    wire N__11352;
    wire N__11347;
    wire N__11346;
    wire N__11345;
    wire N__11344;
    wire N__11341;
    wire N__11336;
    wire N__11331;
    wire N__11326;
    wire N__11325;
    wire N__11324;
    wire N__11323;
    wire N__11322;
    wire N__11321;
    wire N__11318;
    wire N__11313;
    wire N__11306;
    wire N__11299;
    wire N__11296;
    wire N__11293;
    wire N__11290;
    wire N__11287;
    wire N__11284;
    wire N__11281;
    wire N__11278;
    wire N__11275;
    wire N__11272;
    wire N__11269;
    wire N__11268;
    wire N__11267;
    wire N__11266;
    wire N__11259;
    wire N__11256;
    wire N__11251;
    wire N__11248;
    wire N__11245;
    wire N__11242;
    wire N__11239;
    wire N__11236;
    wire N__11233;
    wire N__11230;
    wire N__11227;
    wire N__11224;
    wire N__11221;
    wire N__11218;
    wire N__11215;
    wire N__11212;
    wire N__11209;
    wire N__11206;
    wire N__11203;
    wire N__11200;
    wire N__11197;
    wire N__11196;
    wire N__11191;
    wire N__11188;
    wire N__11185;
    wire N__11184;
    wire N__11179;
    wire N__11176;
    wire N__11175;
    wire N__11172;
    wire N__11169;
    wire N__11166;
    wire N__11161;
    wire N__11160;
    wire N__11155;
    wire N__11152;
    wire N__11151;
    wire N__11146;
    wire N__11143;
    wire N__11140;
    wire N__11139;
    wire N__11136;
    wire N__11135;
    wire N__11132;
    wire N__11127;
    wire N__11122;
    wire N__11121;
    wire N__11120;
    wire N__11119;
    wire N__11114;
    wire N__11109;
    wire N__11104;
    wire N__11101;
    wire N__11098;
    wire N__11095;
    wire N__11092;
    wire N__11089;
    wire N__11086;
    wire N__11083;
    wire N__11080;
    wire N__11077;
    wire N__11076;
    wire N__11073;
    wire N__11070;
    wire N__11065;
    wire N__11064;
    wire N__11061;
    wire N__11058;
    wire N__11055;
    wire N__11050;
    wire N__11047;
    wire N__11046;
    wire N__11043;
    wire N__11040;
    wire N__11035;
    wire N__11032;
    wire N__11029;
    wire N__11028;
    wire N__11027;
    wire N__11024;
    wire N__11023;
    wire N__11022;
    wire N__11011;
    wire N__11008;
    wire N__11005;
    wire N__11002;
    wire N__10999;
    wire N__10996;
    wire N__10993;
    wire N__10990;
    wire N__10987;
    wire N__10984;
    wire N__10981;
    wire N__10978;
    wire N__10975;
    wire N__10974;
    wire N__10969;
    wire N__10966;
    wire N__10965;
    wire N__10964;
    wire N__10957;
    wire N__10954;
    wire N__10951;
    wire N__10948;
    wire N__10945;
    wire N__10942;
    wire N__10939;
    wire N__10936;
    wire N__10933;
    wire N__10930;
    wire \latticehx1k_pll_inst.clk ;
    wire clk_in_c;
    wire GNDG0;
    wire VCCG0;
    wire \uu0.un187_ci_1_cascade_ ;
    wire \uu0.un165_ci_0 ;
    wire \uu0.l_countZ0Z_13 ;
    wire \uu0.l_countZ0Z_12 ;
    wire \uu0.un4_l_count_0_8_cascade_ ;
    wire \uu0.l_countZ0Z_0 ;
    wire \uu0.un44_ci ;
    wire \uu0.un44_ci_cascade_ ;
    wire bfn_1_4_0_;
    wire \buart.Z_tx.un1_bitcount_cry_0 ;
    wire \buart.Z_tx.bitcount_RNIVE1P1_0Z0Z_3 ;
    wire \buart.Z_tx.un1_bitcount_cry_1 ;
    wire \buart.Z_tx.un1_bitcount_cry_2 ;
    wire \buart.Z_tx.bitcount_RNIVE1P1Z0Z_3 ;
    wire \buart.Z_tx.un1_bitcount_axb_3 ;
    wire \buart.Z_tx.un1_bitcount_cry_0_0_c_RNOZ0 ;
    wire \buart.Z_tx.bitcountZ0Z_1 ;
    wire \buart.Z_tx.bitcountZ0Z_3 ;
    wire \buart.Z_tx.bitcountZ0Z_2 ;
    wire \buart.Z_tx.uart_busy_0_i_cascade_ ;
    wire bfn_1_6_0_;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_1 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_2 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_3 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_4 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_5 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_5 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_4 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_6 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_3 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_2 ;
    wire \buart.Z_tx.Z_baudgen.ser_clk_4_cascade_ ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_1 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_0 ;
    wire \Lab_UT.dictrl.N_17_1_cascade_ ;
    wire \Lab_UT.dictrl.g0_i_4_0_cascade_ ;
    wire \Lab_UT.dictrl.N_19 ;
    wire \Lab_UT.dictrl.N_8_2 ;
    wire \Lab_UT.dictrl.N_8_2_cascade_ ;
    wire \Lab_UT.dictrl.g0_i_a8_0_1 ;
    wire \Lab_UT.dictrl.N_1605_1 ;
    wire \Lab_UT.dictrl.currState_0_ret_28_RNOZ0Z_4_cascade_ ;
    wire \Lab_UT.dictrl.N_1605_0 ;
    wire \Lab_UT.dictrl.N_5_0 ;
    wire \Lab_UT.dictrl.g1_0_cascade_ ;
    wire \Lab_UT.dictrl.g0_i_o4_4_1_cascade_ ;
    wire \Lab_UT.dictrl.g0_i_o4_4_cascade_ ;
    wire uart_RXD;
    wire \uu0.l_countZ0Z_2 ;
    wire \uu0.un4_l_count_14_cascade_ ;
    wire \uu0.un4_l_count_13 ;
    wire \uu0.un4_l_count_18_cascade_ ;
    wire \uu0.un4_l_count_0_cascade_ ;
    wire \uu0.un143_ci_0 ;
    wire \uu0.l_countZ0Z_11 ;
    wire \uu0.l_countZ0Z_10 ;
    wire \uu0.un154_ci_9 ;
    wire \uu0.un154_ci_9_cascade_ ;
    wire \uu0.un4_l_count_0_8 ;
    wire \uu0.l_countZ0Z_14 ;
    wire \uu0.l_countZ0Z_8 ;
    wire \uu0.un110_ci ;
    wire \uu0.un198_ci_2 ;
    wire \uu0.un110_ci_cascade_ ;
    wire \uu0.l_countZ0Z_16 ;
    wire \uu0.un220_ci_cascade_ ;
    wire \uu0.l_countZ0Z_9 ;
    wire \uu0.l_countZ0Z_7 ;
    wire \uu0.l_countZ0Z_17 ;
    wire \uu0.l_countZ0Z_3 ;
    wire \uu0.un4_l_count_12 ;
    wire \buart.Z_tx.uart_busy_0_i ;
    wire \buart.Z_tx.ser_clk ;
    wire \buart.Z_tx.bitcountZ0Z_0 ;
    wire \uu0.l_precountZ0Z_2 ;
    wire \uu0.l_precountZ0Z_1 ;
    wire \uu0.l_precountZ0Z_3 ;
    wire \uu0.l_countZ0Z_1 ;
    wire \uu0.l_countZ0Z_18 ;
    wire \uu0.l_countZ0Z_15 ;
    wire \uu0.un4_l_count_11_cascade_ ;
    wire \uu0.un4_l_count_16 ;
    wire \uu2.r_data_wire_0 ;
    wire \uu2.r_data_wire_1 ;
    wire \uu2.r_data_wire_2 ;
    wire \uu2.r_data_wire_3 ;
    wire \uu2.r_data_wire_4 ;
    wire \uu2.r_data_wire_5 ;
    wire \uu2.r_data_wire_6 ;
    wire \uu2.r_data_wire_7 ;
    wire \INVuu2.r_data_reg_0C_net ;
    wire vbuf_tx_data_0;
    wire \buart.Z_tx.shifterZ0Z_1 ;
    wire \buart.Z_tx.shifterZ0Z_0 ;
    wire o_serial_data_c;
    wire vbuf_tx_data_1;
    wire \buart.Z_tx.shifterZ0Z_2 ;
    wire vbuf_tx_data_2;
    wire \buart.Z_tx.shifterZ0Z_3 ;
    wire vbuf_tx_data_3;
    wire \buart.Z_tx.shifterZ0Z_4 ;
    wire vbuf_tx_data_4;
    wire \buart.Z_tx.shifterZ0Z_5 ;
    wire vbuf_tx_data_5;
    wire \buart.Z_tx.shifterZ0Z_6 ;
    wire \INVuu2.vram_rd_clk_det_0C_net ;
    wire \uu2.un1_l_count_1_3_cascade_ ;
    wire \uu2.un1_l_count_1_3 ;
    wire \uu2.un1_l_count_2_0_cascade_ ;
    wire \uu2.l_countZ0Z_2 ;
    wire \uu2.l_countZ0Z_3 ;
    wire \uu2.un306_ci_cascade_ ;
    wire \uu2.un350_ci_cascade_ ;
    wire \uu2.un1_l_count_1_2_0 ;
    wire \uu2.un350_ci ;
    wire \uu2.l_countZ0Z_8 ;
    wire \uu2.l_countZ0Z_5 ;
    wire \uu2.vbuf_count.un328_ci_3 ;
    wire \uu2.vbuf_count.un328_ci_3_cascade_ ;
    wire \uu2.un306_ci ;
    wire \uu2.l_countZ0Z_7 ;
    wire \uu2.l_countZ0Z_6 ;
    wire \uu2.l_countZ0Z_4 ;
    wire \uu2.l_countZ0Z_9 ;
    wire \uu2.un1_l_count_2_2 ;
    wire \Lab_UT.dictrl.N_8_1_cascade_ ;
    wire \Lab_UT.dictrl.N_20_0_cascade_ ;
    wire \Lab_UT.dictrl.N_9_1 ;
    wire \Lab_UT.dictrl.G_30_0_a7_4_1 ;
    wire \Lab_UT.dictrl.G_30_0_a7_1_2 ;
    wire \Lab_UT.dictrl.N_31_0_cascade_ ;
    wire \Lab_UT.dictrl.N_23_1 ;
    wire \Lab_UT.dictrl.G_30_0_2_cascade_ ;
    wire \Lab_UT.dictrl.nextStateZ0Z_1_cascade_ ;
    wire \Lab_UT.dictrl.G_30_0_a7_2_0_cascade_ ;
    wire \Lab_UT.dictrl.G_30_0_0 ;
    wire \Lab_UT.dictrl.G_30_0_a7_0_0 ;
    wire \Lab_UT.dictrl.N_30_0 ;
    wire \Lab_UT.dictrl.i8_mux_0_0_cascade_ ;
    wire \Lab_UT.dictrl.i7_mux_0 ;
    wire \Lab_UT.dictrl.N_12 ;
    wire \Lab_UT.dictrl.G_30_0_a7_2 ;
    wire \Lab_UT.dictrl.N_11_0_cascade_ ;
    wire \Lab_UT.dictrl.N_5_0_0 ;
    wire \Lab_UT.dictrl.g0_4_0_cascade_ ;
    wire \Lab_UT.dictrl.N_8_0_0_cascade_ ;
    wire \Lab_UT.dictrl.N_4 ;
    wire \Lab_UT.dictrl.currState_i_5_2 ;
    wire \Lab_UT.dictrl.G_19_0_a7_4_10_cascade_ ;
    wire \Lab_UT.dictrl.N_21_cascade_ ;
    wire \Lab_UT.dictrl.G_19_0_a7_2_0 ;
    wire \Lab_UT.dictrl.G_19_0_0 ;
    wire \Lab_UT.dictrl.G_19_0_a7_3_2 ;
    wire G_19_0_a7_4_8;
    wire G_19_0_a7_4_1;
    wire \uu0.l_precountZ0Z_0 ;
    wire \uu0.un99_ci_0 ;
    wire \uu0.l_countZ0Z_4 ;
    wire \uu0.l_countZ0Z_5 ;
    wire \uu0.un88_ci_3 ;
    wire \uu0.un66_ci ;
    wire \uu0.un88_ci_3_cascade_ ;
    wire \uu0.l_countZ0Z_6 ;
    wire \uu0.un11_l_count_i_g ;
    wire \uu2.mem0.w_addr_8 ;
    wire \uu2.vram_rd_clk_detZ0Z_1 ;
    wire \uu2.vram_rd_clk_detZ0Z_0 ;
    wire \uu2.vram_rd_clk_det_RNI95711Z0Z_1 ;
    wire \uu2.mem0.w_data_4 ;
    wire \uu2.mem0.w_data_5 ;
    wire \uu2.N_37 ;
    wire \uu2.N_37_cascade_ ;
    wire \uu2.mem0.w_data_3 ;
    wire \uu2.mem0.w_data_1 ;
    wire \uu2.N_51_cascade_ ;
    wire \uu2.N_34 ;
    wire \uu2.N_34_cascade_ ;
    wire \uu2.mem0.w_data_0 ;
    wire \uu2.bitmap_pmux_sn_m15_0_ns_1_cascade_ ;
    wire \uu2.bitmap_pmux_sn_N_65 ;
    wire \uu2.bitmap_pmux_sn_m24_0_ns_1_cascade_ ;
    wire \uu2.bitmap_pmux_sn_i5_mux_cascade_ ;
    wire \uu2.bitmap_pmux_sn_i7_mux_0 ;
    wire \uu2.bitmap_pmux_29_0_cascade_ ;
    wire \uu2.bitmap_pmux ;
    wire \uu2.bitmap_pmux_sn_N_36 ;
    wire vbuf_tx_data_6;
    wire \buart.Z_tx.shifterZ0Z_7 ;
    wire vbuf_tx_data_rdy;
    wire vbuf_tx_data_7;
    wire \buart.Z_tx.shifterZ0Z_8 ;
    wire \buart.Z_tx.un1_uart_wr_i_0_i ;
    wire \uu0.un11_l_count_i ;
    wire \uu2.mem0.w_addr_7 ;
    wire \uu2.mem0.w_addr_1 ;
    wire \uu2.w_data_displaying_2_i_a2_i_a3_1_0 ;
    wire \uu0.un4_l_count_0 ;
    wire \uu2.un1_l_count_2_0 ;
    wire \uu0.delay_lineZ0Z_0 ;
    wire \uu0.delay_lineZ0Z_1 ;
    wire \uu2.l_countZ0Z_1 ;
    wire \uu2.l_countZ0Z_0 ;
    wire \uu2.un284_ci ;
    wire \Lab_UT.dictrl.N_9_cascade_ ;
    wire \Lab_UT.dictrl.N_21_1_cascade_ ;
    wire \Lab_UT.dictrl.g0_0_0_cascade_ ;
    wire \Lab_UT.dictrl.N_1611_0_cascade_ ;
    wire \Lab_UT.dictrl.N_23_0 ;
    wire \Lab_UT.dictrl.N_8_3 ;
    wire \Lab_UT.dictrl.G_28_0_a5_1 ;
    wire \Lab_UT.dictrl.N_19_0 ;
    wire \Lab_UT.dictrl.N_8_3_cascade_ ;
    wire \Lab_UT.dictrl.currState_2_0_rep2_RNIBGCIZ0Z9_cascade_ ;
    wire \Lab_UT.dictrl.G_28_0_0 ;
    wire \Lab_UT.dictrl.currState_2_0_rep2_RNIKH8PZ0Z2 ;
    wire shifter_RNIS6CF1_5;
    wire \Lab_UT.dictrl.m21_rn_1_0_cascade_ ;
    wire \Lab_UT.dictrl.m21_rn_0 ;
    wire \Lab_UT.dictrl.g1_0_1 ;
    wire \Lab_UT.dictrl.N_7_1 ;
    wire \Lab_UT.dictrl.nextState_0_1 ;
    wire \Lab_UT.dictrl.N_20_cascade_ ;
    wire \Lab_UT.dictrl.decoder.g0Z0Z_5_cascade_ ;
    wire \Lab_UT.dictrl.decoder.g0Z0Z_1 ;
    wire \Lab_UT.dictrl.N_36_1_cascade_ ;
    wire G_28_0_a5_0_4_cascade_;
    wire shifter_RNI1D8L1_4;
    wire bfn_4_16_0_;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_1 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_2 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_3 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_4 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_5 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_2 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_1 ;
    wire \uu2.trig_rd_is_det_cascade_ ;
    wire \uu2.trig_rd_detZ0Z_1 ;
    wire \uu2.vram_rd_clkZ0 ;
    wire \uu2.un1_l_count_1_0 ;
    wire \uu2.trig_rd_detZ0Z_0 ;
    wire \uu2.vbuf_raddr.un448_ci_0 ;
    wire \uu2.vbuf_raddr.un426_ci_3_cascade_ ;
    wire \uu2.r_addrZ0Z_8 ;
    wire \uu2.vbuf_raddr.un426_ci_3 ;
    wire \uu2.r_addrZ0Z_7 ;
    wire \uu2.un404_ci_0_cascade_ ;
    wire \uu2.r_addrZ0Z_6 ;
    wire \uu2.r_addrZ0Z_2 ;
    wire \uu2.r_addrZ0Z_1 ;
    wire \uu2.r_addrZ0Z_0 ;
    wire \uu2.r_addrZ0Z_3 ;
    wire \uu2.trig_rd_is_det_0 ;
    wire \uu2.bitmap_pmux_sn_N_42 ;
    wire \uu2.bitmap_pmux_26_bm_1_cascade_ ;
    wire \uu2.N_161 ;
    wire \uu2.N_400_cascade_ ;
    wire \uu2.N_409 ;
    wire \uu2.bitmap_RNI1PH82Z0Z_34 ;
    wire \uu2.N_404 ;
    wire \uu2.bitmapZ0Z_290 ;
    wire \uu2.bitmapZ0Z_40 ;
    wire \uu2.bitmapZ0Z_296 ;
    wire \INVuu2.bitmap_290C_net ;
    wire \uu2.bitmap_pmux_25_am_1_cascade_ ;
    wire \uu2.bitmapZ0Z_197 ;
    wire \uu2.bitmapZ0Z_66 ;
    wire \INVuu2.bitmap_197C_net ;
    wire \uu2.bitmap_RNI2JA82Z0Z_212_cascade_ ;
    wire \uu2.N_31_i ;
    wire \uu2.bitmap_RNIM7D32Z0Z_69 ;
    wire \uu2.bitmap_pmux_27_ns_1_cascade_ ;
    wire \uu2.N_407 ;
    wire \Lab_UT.segmentUQ_0_0_cascade_ ;
    wire \Lab_UT.N_65_0_cascade_ ;
    wire \Lab_UT.segment_1_0_6 ;
    wire \Lab_UT.N_76_0_cascade_ ;
    wire \INVuu2.bitmap_72C_net ;
    wire \uu2.bitmapZ0Z_72 ;
    wire \uu2.bitmapZ0Z_200 ;
    wire \uu2.bitmap_RNIOS152Z0Z_72 ;
    wire \Lab_UT.dictrl.currState_ret_RNI7FNUZ0 ;
    wire \Lab_UT.Mone_at_0_cascade_ ;
    wire \Lab_UT.N_77_0 ;
    wire \Lab_UT.dictrl.N_23 ;
    wire \Lab_UT.dictrl.N_23_cascade_ ;
    wire \Lab_UT.dictrl.nextState_RNIA8EV3Z0Z_1 ;
    wire \Lab_UT.dictrl.N_10 ;
    wire \Lab_UT.dictrl.N_12_0_cascade_ ;
    wire \Lab_UT.dictrl.G_28_0_a5_2_1 ;
    wire \Lab_UT.dictrl.dicLdAMtensZ0 ;
    wire \Lab_UT.dictrl.dicLdAMtens_rst ;
    wire \Lab_UT.dictrl.r_dicLdMtens16_1 ;
    wire \Lab_UT.dictrl.g0_10_0_N_4L6_1_cascade_ ;
    wire \Lab_UT.dictrl.r_dicLdMtens17_1 ;
    wire \Lab_UT.dictrl.r_dicLdMtens22_2 ;
    wire \Lab_UT.dictrl.N_34_cascade_ ;
    wire \Lab_UT.dictrl.currState_2_RNI0P25DZ0Z_1 ;
    wire \Lab_UT.dictrl.m15_bm_cascade_ ;
    wire \Lab_UT.dictrl.nextState_0_0 ;
    wire \Lab_UT.dictrl.N_7_0 ;
    wire \Lab_UT.dictrl.N_1609_1 ;
    wire \Lab_UT.dictrl.N_38 ;
    wire \Lab_UT.dictrl.currState_ret_5_RNOZ0Z_0 ;
    wire \Lab_UT.dictrl.N_23_0_0 ;
    wire \Lab_UT.dictrl.N_13_0_0 ;
    wire \Lab_UT.dictrl.N_14_0_0_0_cascade_ ;
    wire \Lab_UT.dictrl.N_1609_0_0 ;
    wire \Lab_UT.dictrl.N_8 ;
    wire \Lab_UT.dictrl.N_7 ;
    wire \Lab_UT.dictrl.N_9_0_cascade_ ;
    wire \Lab_UT.dictrl.g0_6 ;
    wire \Lab_UT.dictrl.N_6_0 ;
    wire \Lab_UT.dictrl.N_9 ;
    wire \Lab_UT.dictrl.m15_am ;
    wire \Lab_UT.dictrl.N_20_1 ;
    wire \Lab_UT.dictrl.currState_0_rep1 ;
    wire \buart.Z_rx.bitcount_fast_es_RNIAJ1GZ0Z_3_cascade_ ;
    wire bu_rx_data_rdy_cascade_;
    wire \Lab_UT.dictrl.N_5_0_1 ;
    wire \Lab_UT.dictrl.g0_3_1_cascade_ ;
    wire \Lab_UT.dictrl.g0_1_0_0 ;
    wire bu_rx_data_fast_0;
    wire \Lab_UT.dictrl.de_num_1_2 ;
    wire bu_rx_data_fast_7;
    wire \Lab_UT.dictrl.decoder.g0_5_0_cascade_ ;
    wire \Lab_UT.dictrl.de_cr_0_0 ;
    wire \Lab_UT.dictrl.decoder.g0_6_0 ;
    wire bu_rx_data_fast_6;
    wire \Lab_UT.dictrl.decoder.g0Z0Z_4 ;
    wire bu_rx_data_fast_4;
    wire bu_rx_data_fast_5;
    wire \buart.Z_rx.hhZ0Z_0 ;
    wire \Lab_UT.dictrl.decoder.g0Z0Z_7_cascade_ ;
    wire \Lab_UT.dictrl.currState_fast_0 ;
    wire \Lab_UT.dictrl.g1_4_1_0_cascade_ ;
    wire \Lab_UT.dictrl.de_littleA_0 ;
    wire \Lab_UT.dictrl.g1_4_cascade_ ;
    wire \Lab_UT.dictrl.N_17_0_0 ;
    wire \Lab_UT.dictrl.decoder.g0_5_1 ;
    wire \Lab_UT.dictrl.m7_sx ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_3 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_0 ;
    wire \buart.Z_rx.Z_baudgen.ser_clk_3 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO ;
    wire \buart.Z_rx.ser_clk_cascade_ ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_4 ;
    wire \resetGen.reset_count_2_0_4_cascade_ ;
    wire \uu2.mem0.w_addr_2 ;
    wire \uu2.mem0.w_addr_4 ;
    wire \uu2.mem0.w_addr_5 ;
    wire \uu2.mem0.w_addr_6 ;
    wire \uu2.bitmap_pmux_sn_N_20 ;
    wire \uu2.bitmapZ0Z_168 ;
    wire \uu2.N_17_cascade_ ;
    wire \uu2.bitmap_RNIELSJ2Z0Z_111 ;
    wire \uu2.bitmap_pmux_sn_N_54_mux ;
    wire \uu2.bitmapZ0Z_111 ;
    wire \INVuu2.bitmap_111C_net ;
    wire \uu2.bitmap_pmux_sn_N_33 ;
    wire \uu2.N_39_cascade_ ;
    wire \uu2.N_48 ;
    wire \INVuu2.w_addr_displaying_nesr_3C_net ;
    wire \uu2.bitmap_pmux_24_am_1 ;
    wire \uu2.bitmapZ0Z_87 ;
    wire \uu2.N_386_cascade_ ;
    wire \uu2.w_addr_displaying_nesr_RNI1JET2Z0Z_7_cascade_ ;
    wire \uu2.bitmapZ0Z_314 ;
    wire \uu2.bitmap_pmux_23_ns_1 ;
    wire \uu2.bitmap_pmux_sn_N_15 ;
    wire \uu2.w_addr_displayingZ0Z_2 ;
    wire \INVuu2.bitmap_87C_net ;
    wire \Lab_UT.L3_segment3_0_i_1_0 ;
    wire \Lab_UT.L3_segment3_0_i_1_3 ;
    wire \Lab_UT.L3_segment3_1_2_cascade_ ;
    wire \Lab_UT.Mone_at_0 ;
    wire \Lab_UT.Mone_at_3 ;
    wire \Lab_UT.Mone_at_2 ;
    wire \Lab_UT.Mone_at_1 ;
    wire \Lab_UT.L3_segment3_1_1_cascade_ ;
    wire \uu2.bitmapZ0Z_203 ;
    wire \uu2.bitmapZ0Z_75 ;
    wire \uu2.bitmap_pmux_24_bm_1 ;
    wire \INVuu2.bitmap_203C_net ;
    wire \Lab_UT.N_76_cascade_ ;
    wire \uu2.bitmapZ0Z_194 ;
    wire \Lab_UT.L3_segment4_1_1_cascade_ ;
    wire \uu2.bitmapZ0Z_69 ;
    wire \Lab_UT.L3_segment4_1_0 ;
    wire \uu2.bitmapZ0Z_34 ;
    wire \Lab_UT.segment_1_6_cascade_ ;
    wire \uu2.bitmapZ0Z_162 ;
    wire \INVuu2.bitmap_194C_net ;
    wire \Lab_UT.dictrl.N_1614_0 ;
    wire \Lab_UT.dictrl.N_26 ;
    wire \Lab_UT.dictrl.un1_currState_6 ;
    wire \Lab_UT.dictrl.r_enableZ0Z1 ;
    wire \Lab_UT.dictrl.enableSeg3 ;
    wire \Lab_UT.dictrl.r_enableZ0Z3 ;
    wire \Lab_UT.dictrl.enableSeg4 ;
    wire \Lab_UT.dictrl.un1_currState_7 ;
    wire \Lab_UT.dictrl.r_enableZ0Z4 ;
    wire \Lab_UT.dictrl.N_1605_1_0 ;
    wire \Lab_UT.dictrl.N_36_0_cascade_ ;
    wire \Lab_UT.dictrl.nextStateZ0Z_3_cascade_ ;
    wire \Lab_UT.dictrl.r_dicLdMtens21_1 ;
    wire \Lab_UT.dictrl.N_18 ;
    wire \Lab_UT.dictrl.N_33 ;
    wire \Lab_UT.dictrl.N_1607_0_0 ;
    wire \Lab_UT.dictrl.N_10_0_0 ;
    wire \Lab_UT.dictrl.g1 ;
    wire \Lab_UT.dictrl.g2_cascade_ ;
    wire \Lab_UT.dictrl.nextState_RNO_9Z0Z_1_cascade_ ;
    wire \Lab_UT.dictrl.g0_i_a4_1 ;
    wire \Lab_UT.dictrl.nextState_RNO_4Z0Z_1_cascade_ ;
    wire \Lab_UT.dictrl.nextState_RNO_3Z0Z_1 ;
    wire \Lab_UT.dictrl.g0_i_o4_5 ;
    wire \Lab_UT.dictrl.N_11 ;
    wire \Lab_UT.dictrl.N_18_0 ;
    wire \Lab_UT.dictrl.g1_3_0 ;
    wire \Lab_UT.dictrl.N_13_0 ;
    wire \Lab_UT.dictrl.g1_4_0_cascade_ ;
    wire \Lab_UT.dictrl.N_14 ;
    wire \Lab_UT.dictrl.r_dicLdMtens20_0_cascade_ ;
    wire \Lab_UT.dictrl.N_6ctr ;
    wire \Lab_UT.dictrl.r_dicLdMtens22_2_reti ;
    wire \Lab_UT.dictrl.N_7_1_0 ;
    wire \Lab_UT.dictrl.r_dicLdMtens22_2_reti_cascade_ ;
    wire \Lab_UT.dictrl.g0_0_3 ;
    wire \Lab_UT.dictrl.N_10ctr ;
    wire \Lab_UT.dictrl.r_dicLdMtens22_4_0 ;
    wire N_7;
    wire \Lab_UT.dictrl.N_20 ;
    wire \Lab_UT.dictrl.de_littleA ;
    wire Lab_UT_dictrl_decoder_de_cr_1_cascade_;
    wire \Lab_UT.dictrl.N_30 ;
    wire \Lab_UT.dictrl.N_41_mux ;
    wire \Lab_UT.dictrl.N_34 ;
    wire \Lab_UT.dictrl.N_31_cascade_ ;
    wire \Lab_UT.dictrl.nextState_0_2 ;
    wire \Lab_UT.dictrl.currState_0_ret_29_RNIDFRSEEZ0 ;
    wire buart__rx_bitcount_fast_2;
    wire buart__rx_bitcount_fast_4;
    wire buart__rx_bitcount_fast_3;
    wire \Lab_UT.dictrl.decoder.g0_6_1 ;
    wire \buart.Z_rx.un1_sample_0_cascade_ ;
    wire \buart.Z_rx.sample ;
    wire \buart.Z_rx.idle_0_cascade_ ;
    wire \buart.Z_rx.idle ;
    wire \buart.Z_rx.ser_clk ;
    wire \buart.Z_rx.idle_cascade_ ;
    wire \buart.Z_rx.N_27_0_i ;
    wire \buart.Z_rx.startbit ;
    wire \buart.Z_rx.bitcounte_0_0 ;
    wire buart__rx_bitcount_0;
    wire bfn_6_16_0_;
    wire buart__rx_bitcount_1;
    wire \buart.Z_rx.bitcount_cry_0_THRU_CO ;
    wire \buart.Z_rx.bitcount_cry_0 ;
    wire \buart.Z_rx.bitcount_cry_1_THRU_CO ;
    wire \buart.Z_rx.bitcount_cry_1 ;
    wire \buart.Z_rx.bitcount_cry_2_THRU_CO ;
    wire \buart.Z_rx.bitcount_cry_2 ;
    wire \buart.Z_rx.bitcount_cry_3 ;
    wire \buart.Z_rx.bitcount_cry_3_THRU_CO ;
    wire \Lab_UT.uu0.l_countZ0Z_13 ;
    wire \Lab_UT.uu0.un143_ci_0_cascade_ ;
    wire \Lab_UT.uu0.un154_ci_9_cascade_ ;
    wire \Lab_UT.uu0.l_countZ0Z_12 ;
    wire \Lab_UT.uu0.un165_ci_0 ;
    wire \uu2.un3_w_addr_user_4_cascade_ ;
    wire \uu2.un3_w_addr_user_5 ;
    wire \uu2.w_addr_displayingZ0Z_3 ;
    wire \uu2.mem0.w_addr_3 ;
    wire \uu2.vbuf_w_addr_user.un448_ci_0_cascade_ ;
    wire \uu2.w_addr_userZ0Z_8 ;
    wire \uu2.w_addr_userZ0Z_7 ;
    wire \INVuu2.w_addr_user_nesr_3C_net ;
    wire \uu2.w_addr_displayingZ0Z_1 ;
    wire \uu2.N_39 ;
    wire \INVuu2.w_addr_displaying_8C_net ;
    wire \uu2.w_addr_displayingZ0Z_5 ;
    wire \uu2.w_addr_displayingZ0Z_4 ;
    wire \uu2.N_41 ;
    wire \uu2.w_addr_displayingZ0Z_6 ;
    wire \uu2.N_41_cascade_ ;
    wire \uu2.N_43 ;
    wire \uu2.N_40 ;
    wire \uu2.N_43_cascade_ ;
    wire \uu2.w_addr_displaying_RNIFCPV4Z0Z_8 ;
    wire \uu2.w_addr_displaying_RNIFCPV4Z0Z_8_cascade_ ;
    wire \uu2.N_36_0 ;
    wire \Lab_UT.L3_segment2_1_1 ;
    wire \Lab_UT.L3_segment2_0_i_1_3_cascade_ ;
    wire \Lab_UT.L3_segment2_1_2_cascade_ ;
    wire \uu2.bitmapZ0Z_215 ;
    wire \Lab_UT.L3_segment2_0_i_1_0_cascade_ ;
    wire \INVuu2.bitmap_308C_net ;
    wire \uu2.bitmapZ0Z_52 ;
    wire \uu2.w_addr_displayingZ0Z_8 ;
    wire \uu2.bitmapZ0Z_308 ;
    wire \uu2.N_158 ;
    wire \Lab_UT.segmentUQ_0_0_1_cascade_ ;
    wire \Lab_UT.N_65_2_cascade_ ;
    wire \Lab_UT.segment_1_2_6 ;
    wire \uu2.bitmapZ0Z_186 ;
    wire \Lab_UT.N_76_2_cascade_ ;
    wire \INVuu2.bitmap_90C_net ;
    wire \uu2.bitmapZ0Z_90 ;
    wire \uu2.bitmapZ0Z_218 ;
    wire \uu2.w_addr_displayingZ0Z_7 ;
    wire \Lab_UT.N_76_1_cascade_ ;
    wire \uu2.bitmapZ0Z_212 ;
    wire \Lab_UT.N_65_1_cascade_ ;
    wire \Lab_UT.segment_1_1_6 ;
    wire \uu2.bitmapZ0Z_180 ;
    wire \Lab_UT.N_77_1 ;
    wire \uu2.bitmapZ0Z_84 ;
    wire \INVuu2.bitmap_212C_net ;
    wire \Lab_UT.L3_segment4_0_i_1_5 ;
    wire \Lab_UT.N_65 ;
    wire \Lab_UT.Mten_at_3_cascade_ ;
    wire \Lab_UT.segment_1_3 ;
    wire \Lab_UT.N_69_0 ;
    wire \Lab_UT.N_69_0_cascade_ ;
    wire \Lab_UT.N_92 ;
    wire \Lab_UT.N_67_0 ;
    wire \Lab_UT.N_91 ;
    wire \Lab_UT.N_83 ;
    wire \Lab_UT.Mten_at_0 ;
    wire \Lab_UT.Mten_at_3 ;
    wire \Lab_UT.Mten_at_0_cascade_ ;
    wire \Lab_UT.N_77 ;
    wire \Lab_UT.Mten_at_1 ;
    wire \Lab_UT.dictrl.g0_13_1 ;
    wire \Lab_UT.dictrl.g0_1 ;
    wire \Lab_UT.dictrl.g0_i_o4_0_0 ;
    wire \Lab_UT.dictrl.currState_0_ret_20and_1_0_cascade_ ;
    wire \Lab_UT.dictrl.de_cr ;
    wire \Lab_UT.dictrl.N_13 ;
    wire \Lab_UT.dictrl.N_17_0 ;
    wire \Lab_UT.dictrl.N_13_cascade_ ;
    wire \Lab_UT.dictrl.G_19_0_2 ;
    wire \Lab_UT.dictrl.nextStateZ0Z_2_cascade_ ;
    wire \Lab_UT.dictrl.dicLdASones_rst ;
    wire \Lab_UT.dictrl.dicLdASones_rst_cascade_ ;
    wire \Lab_UT.dictrl.dicLdASonesZ0 ;
    wire \Lab_UT.dictrl.N_5ctr ;
    wire \Lab_UT.dictrl.N_7ctr ;
    wire \Lab_UT.dictrl.nextState_RNIGHD18Z0Z_1 ;
    wire \Lab_UT.dictrl.i8_mux ;
    wire \Lab_UT.dictrl.currState_2_RNI1O2A_0Z0Z_1 ;
    wire \Lab_UT.dictrl.r_dicLdMtens15_1i_cascade_ ;
    wire \Lab_UT.dictrl.currState_ret_3and ;
    wire \Lab_UT.dictrl.currState_0_ret_28_RNOZ0Z_2 ;
    wire \Lab_UT.dictrl.N_8ctr ;
    wire \Lab_UT.dictrl.currState_0_ret_28_RNOZ0Z_3_cascade_ ;
    wire \Lab_UT.dictrl.N_8_0 ;
    wire \Lab_UT.dictrl.r_dicLdMtens21_1_reti ;
    wire \Lab_UT.dictrl.decoder.de_littleA_2Z0Z_0 ;
    wire \Lab_UT.dictrl.de_littleA_1_cascade_ ;
    wire \Lab_UT.dictrl.N_37_0_cascade_ ;
    wire \Lab_UT.dictrl.g0_15_rn_1 ;
    wire \Lab_UT.dictrl.G_19_0_a7_0_1 ;
    wire G_19_0_a7_4_7;
    wire \Lab_UT.dictrl.currState_2_RNIEPCJZ0Z_1 ;
    wire \Lab_UT.dictrl.nextState_0_3 ;
    wire \Lab_UT.dictrl.N_1612_0 ;
    wire \Lab_UT.dictrl.currState_2_RNI2P2AZ0Z_2 ;
    wire Lab_UT_dictrl_currState_1;
    wire \Lab_UT.dictrl.G_19_0_a7_2 ;
    wire \Lab_UT.dictrl.decoder.g0_2Z0Z_2 ;
    wire Lab_UT_dictrl_decoder_de_cr_2_cascade_;
    wire buart__rx_bitcount_2_rep1;
    wire \Lab_UT.dictrl.decoder.g0_4_0_cascade_ ;
    wire \Lab_UT.dictrl.de_cr_1_0 ;
    wire \Lab_UT.dictrl.de_cr_0 ;
    wire bu_rx_data_fast_2;
    wire \Lab_UT.dictrl.decoder.g0_3Z0Z_0 ;
    wire \Lab_UT.dictrl.de_cr_1_2 ;
    wire \Lab_UT.dictrl.decoder.g0_4Z0Z_3 ;
    wire \Lab_UT.dictrl.decoder.g0_3_2_cascade_ ;
    wire Lab_UT_dictrl_decoder_de_cr_1_1;
    wire \Lab_UT.dictrl.de_cr_2_0 ;
    wire \Lab_UT.dictrl.decoder.g0_4_1 ;
    wire buart__rx_bitcount_4;
    wire buart__rx_bitcount_3;
    wire buart__rx_bitcount_2;
    wire \Lab_UT.dictrl.g0_8_cascade_ ;
    wire buart__rx_valid_2_0;
    wire \Lab_UT.dictrl.g0_11 ;
    wire \Lab_UT.uu0.un99_ci_0_cascade_ ;
    wire \Lab_UT.uu0.un88_ci_3 ;
    wire \Lab_UT.uu0.un88_ci_3_cascade_ ;
    wire \Lab_UT.uu0.l_countZ0Z_7 ;
    wire \Lab_UT.uu0.l_countZ0Z_17 ;
    wire \Lab_UT.uu0.un110_ci_cascade_ ;
    wire \Lab_UT.uu0.un220_ci ;
    wire \Lab_UT.uu0.l_countZ0Z_9 ;
    wire \Lab_UT.uu0.l_countZ0Z_10 ;
    wire \Lab_UT.uu0.un4_l_count_14_cascade_ ;
    wire \Lab_UT.uu0.un187_ci_1_cascade_ ;
    wire \Lab_UT.uu0.un154_ci_9 ;
    wire \Lab_UT.uu0.l_countZ0Z_14 ;
    wire \Lab_UT.uu0.un4_l_count_0_8 ;
    wire \Lab_UT.uu0.un198_ci_2 ;
    wire \Lab_UT.uu0.un110_ci ;
    wire \Lab_UT.uu0.l_countZ0Z_8 ;
    wire \uu2.un28_w_addr_user_i_0 ;
    wire \uu2.un1_w_user_lf_0_cascade_ ;
    wire \uu2.vram_wr_en_0_iZ0 ;
    wire \uu2.un1_w_user_lf_0 ;
    wire \uu2.un3_w_addr_user ;
    wire \uu2.un1_w_user_cr_0 ;
    wire \uu2.un1_w_user_cr_0_cascade_ ;
    wire \uu2.N_71 ;
    wire \uu2.un4_w_user_data_rdyZ0Z_0_cascade_ ;
    wire \uu2.mem0.w_data_6 ;
    wire \uu2.un1_w_user_crZ0Z_4 ;
    wire \uu2.un1_w_user_lfZ0Z_4 ;
    wire \uu2.mem0.w_data_2 ;
    wire \uu2.un4_w_user_data_rdyZ0Z_0 ;
    wire \uu2.mem0.w_addr_0 ;
    wire \INVuu2.w_addr_user_0C_net ;
    wire \uu2.w_addr_userZ0Z_0 ;
    wire \uu2.w_addr_userZ0Z_2 ;
    wire \uu2.w_addr_userZ0Z_3 ;
    wire \uu2.w_addr_userZ0Z_1 ;
    wire \resetGen.un252_ci_cascade_ ;
    wire \resetGen.reset_countZ0Z_3 ;
    wire \resetGen.reset_countZ0Z_1 ;
    wire \resetGen.reset_countZ0Z_0 ;
    wire \resetGen.un241_ci ;
    wire \resetGen.reset_countZ0Z_4 ;
    wire \resetGen.un241_ci_cascade_ ;
    wire \resetGen.reset_countZ0Z_2 ;
    wire \Lab_UT.uu0.delay_lineZ0Z_1 ;
    wire \Lab_UT.uu0.un11_l_count_i ;
    wire \Lab_UT.L3_segment1_1_0_3 ;
    wire \Lab_UT.L3_segment1_0_i_1_0_cascade_ ;
    wire \uu2.bitmapZ0Z_58 ;
    wire \Lab_UT.L3_segment1_0_i_1_1 ;
    wire \Lab_UT.dictrl.enableSeg1 ;
    wire \Lab_UT.L3_segment1_1_2_cascade_ ;
    wire \INVuu2.bitmap_93C_net ;
    wire \uu2.bitmapZ0Z_93 ;
    wire \uu2.bitmap_pmux_25_bm_1 ;
    wire \uu2.bitmapZ0Z_221 ;
    wire \uu2.w_addr_displayingZ0Z_0 ;
    wire \uu2.bitmap_RNI1D952Z0Z_93 ;
    wire \Lab_UT.Sone_at_0 ;
    wire \Lab_UT.Sone_at_0_cascade_ ;
    wire \Lab_UT.N_77_2 ;
    wire \Lab_UT.Sone_at_3 ;
    wire \Lab_UT.Sone_at_2 ;
    wire \Lab_UT.Sten_at_1 ;
    wire \Lab_UT.Sten_at_0 ;
    wire \Lab_UT.Sten_at_3 ;
    wire \Lab_UT.Sten_at_1_cascade_ ;
    wire \Lab_UT.Sten_at_2 ;
    wire \Lab_UT.segmentUQ_0_0_0 ;
    wire \Lab_UT.dictrl.L3_segment1_1 ;
    wire \Lab_UT.Sone_at_1 ;
    wire \Lab_UT.dictrl.r_enable1_2_i_m ;
    wire \Lab_UT.alarm_or_time_0 ;
    wire \Lab_UT.alarm_or_time_0_cascade_ ;
    wire \Lab_UT.Mten_at_2 ;
    wire \Lab_UT.dictrl.r_enable1_2_m ;
    wire \Lab_UT.dictrl.r_enable1_2_m_cascade_ ;
    wire \Lab_UT.dictrl.g0_i_a4_0 ;
    wire \Lab_UT.dictrl.r_enableZ0Z2 ;
    wire \Lab_UT.dictrl.enableSeg2 ;
    wire \Lab_UT.dictrl.currState_0_ret_20and_1_0 ;
    wire \Lab_UT.dictrl.r_dicLdMtens16_reti ;
    wire \Lab_UT.dictrl.r_dicLdMtens19 ;
    wire \Lab_UT.dictrl.r_dicLdMtens22_i_6 ;
    wire \Lab_UT.dictrl.r_enable2_3_iv_0_cascade_ ;
    wire \Lab_UT.dictrl.r_enable2_3_iv_3 ;
    wire \Lab_UT.dictrl.r_Sone_init17_4 ;
    wire \Lab_UT.dictrl.r_dicLdMtens23_i_6 ;
    wire \Lab_UT.dictrl.un1_r_dicLdMtens19_0_cascade_ ;
    wire \Lab_UT.dictrl.r_alarm_or_timeZ0 ;
    wire \Lab_UT.dictrl.r_dicLdMtens18_i_6 ;
    wire \Lab_UT.dictrl.r_dicLdMtens17_i_6 ;
    wire \Lab_UT.dictrl.r_dicLdMtens16 ;
    wire \Lab_UT.dictrl.nextStateZ0Z_2 ;
    wire \Lab_UT.dictrl.nextStateZ0Z_1 ;
    wire \Lab_UT.dictrl.r_dicLdMtens17 ;
    wire \Lab_UT.dictrl.currState_ret_1and ;
    wire \Lab_UT.dictrl.dicLdAMones_rst ;
    wire \Lab_UT.dictrl.dicLdAMonesZ0 ;
    wire \Lab_UT.dictrl.dicLdAMones_rst_cascade_ ;
    wire \Lab_UT.dictrl.r_dicLdMtens23_2 ;
    wire \Lab_UT.dictrl.dicLdAStensZ0 ;
    wire \Lab_UT.dictrl.dicLdAStens_rst ;
    wire \resetGen.escKeyZ0 ;
    wire \Lab_UT.dictrl.currState_3_rep1 ;
    wire \Lab_UT.dictrl.N_5 ;
    wire \Lab_UT.dictrl.N_6 ;
    wire \Lab_UT.dictrl.r_dicLdMtens14_i_6 ;
    wire \Lab_UT.dictrl.r_dicLdMtens20_i_6 ;
    wire \Lab_UT.dictrl.r_enable3_3_iv_1 ;
    wire \buart.Z_rx.G_30_0_o3_1_0_cascade_ ;
    wire Lab_UT_dictrl_decoder_de_cr_1;
    wire \Lab_UT.dictrl.currStateZ0Z_0 ;
    wire N_6_cascade_;
    wire \Lab_UT.dictrl.N_21_0 ;
    wire \resetGen.escKey_4_0 ;
    wire \Lab_UT.dictrl.nextStateZ0Z_0 ;
    wire \Lab_UT.dictrl.currState_0_rep2 ;
    wire \Lab_UT.dictrl.g0_7_cascade_ ;
    wire \Lab_UT.dictrl.g0_10 ;
    wire bu_rx_data_fast_1;
    wire bu_rx_data_3_rep1;
    wire \Lab_UT.dictrl.g1_5_1_cascade_ ;
    wire \Lab_UT.dictrl.g1_7_1 ;
    wire bu_rx_data_2_rep1;
    wire \Lab_UT.dictrl.g1_4_1 ;
    wire \Lab_UT.dictrl.currState_fast_3 ;
    wire \buart.Z_rx.G_30_0_o3_1_4 ;
    wire \Lab_UT.dictrl.nextStateZ0Z_3 ;
    wire bu_rx_data_4_rep1;
    wire bu_rx_data_1_rep1;
    wire \Lab_UT.dictrl.decoder.g0Z0Z_3 ;
    wire bu_rx_data_0_rep1;
    wire bu_rx_data_6_rep1;
    wire bu_rx_data_5_rep1;
    wire bu_rx_data_fast_3;
    wire \buart.Z_rx.hhZ0Z_1 ;
    wire bu_rx_data_7_rep1;
    wire \Lab_UT.uu0.un44_ci ;
    wire \Lab_UT.uu0.un44_ci_cascade_ ;
    wire \Lab_UT.uu0.l_countZ0Z_3 ;
    wire \Lab_UT.uu0.l_countZ0Z_2 ;
    wire \Lab_UT.uu0.un66_ci_cascade_ ;
    wire \Lab_UT.uu0.l_countZ0Z_4 ;
    wire \Lab_UT.uu0.un66_ci ;
    wire \Lab_UT.uu0.un11_l_count_i_g ;
    wire \Lab_UT.uu0.delay_lineZ0Z_0 ;
    wire \Lab_UT.uu0.l_countZ0Z_5 ;
    wire \Lab_UT.uu0.l_precountZ0Z_3 ;
    wire \Lab_UT.uu0.l_countZ0Z_1 ;
    wire \Lab_UT.uu0.l_countZ0Z_18 ;
    wire \Lab_UT.uu0.l_countZ0Z_15 ;
    wire \Lab_UT.uu0.un4_l_count_11_cascade_ ;
    wire \Lab_UT.uu0.l_countZ0Z_6 ;
    wire \Lab_UT.uu0.un4_l_count_12 ;
    wire \Lab_UT.uu0.un4_l_count_16_cascade_ ;
    wire \Lab_UT.uu0.un4_l_count_18 ;
    wire \Lab_UT.uu0.l_precountZ0Z_1 ;
    wire \Lab_UT.uu0.l_countZ0Z_16 ;
    wire \Lab_UT.uu0.l_countZ0Z_11 ;
    wire \Lab_UT.uu0.l_precountZ0Z_2 ;
    wire \Lab_UT.uu0.l_countZ0Z_0 ;
    wire \Lab_UT.uu0.un4_l_count_13 ;
    wire \uu2.w_addr_userZ0Z_5 ;
    wire \uu2.w_addr_userZ0Z_4 ;
    wire \uu2.un28_w_addr_user_i ;
    wire \uu2.un404_ci ;
    wire \uu2.un426_ci_3 ;
    wire \uu2.w_addr_userZ0Z_6 ;
    wire \INVuu2.w_addr_user_5C_net ;
    wire \uu2.w_addr_user_RNIMJ3O2Z0Z_2 ;
    wire L3_tx_data_rdy;
    wire L3_tx_data_6;
    wire \Lab_UT.display.N_88_cascade_ ;
    wire L3_tx_data_1;
    wire \Lab_UT.display.N_120_cascade_ ;
    wire L3_tx_data_4;
    wire L3_tx_data_5;
    wire \Lab_UT.display.N_153_cascade_ ;
    wire \Lab_UT.display.dOutP_0_iv_i_1_1 ;
    wire \Lab_UT.display.N_150 ;
    wire \Lab_UT.display.N_101_cascade_ ;
    wire \Lab_UT.display.N_88 ;
    wire \Lab_UT.display.dOutP_0_iv_i_0_3_cascade_ ;
    wire \Lab_UT.display.dOutP_0_iv_i_2_3 ;
    wire L3_tx_data_3;
    wire \uu2.r_addrZ0Z_5 ;
    wire \Lab_UT.di_AMones_0 ;
    wire \Lab_UT.di_AMones_2 ;
    wire \Lab_UT.ld_enable_AMones ;
    wire \Lab_UT.di_AMones_3 ;
    wire \Lab_UT.di_ASones_0 ;
    wire \Lab_UT.di_ASones_1 ;
    wire \Lab_UT.di_ASones_2 ;
    wire \Lab_UT.ld_enable_AMtens ;
    wire \Lab_UT.di_AStens_3 ;
    wire \Lab_UT.ld_enable_ASones ;
    wire \Lab_UT.di_ASones_3 ;
    wire \Lab_UT.ld_enable_AStens ;
    wire \Lab_UT.uu0.un4_l_count_0 ;
    wire \Lab_UT.halfPulse ;
    wire \Lab_UT.displayAlarmZ0Z_1 ;
    wire \Lab_UT.dicLdStens ;
    wire \Lab_UT.dicLdStens_latmux ;
    wire \Lab_UT.didp.Stens_subtractor.un1_q_axb0 ;
    wire \Lab_UT.didp.Stens_subtractor.q_RNO_0_0_3 ;
    wire \Lab_UT.didp.Stens_subtractor.N_86 ;
    wire \Lab_UT.didp.Stens_subtractor.q_RNO_0_1_2 ;
    wire \Lab_UT.didp.q_RNIDDF11_3_cascade_ ;
    wire led_c_3;
    wire \Lab_UT.didp.q_RNI1TVP_3 ;
    wire \Lab_UT.didp.q_RNIBBF11_2 ;
    wire \Lab_UT.didp.q_RNIVQVP_2 ;
    wire led_c_2;
    wire \Lab_UT.dictrl.r_Sone_init5 ;
    wire Lab_UT_dictrl_r_Sone_init17;
    wire \Lab_UT.dictrl.r_dicAlarmTrigZ0 ;
    wire \Lab_UT.displayAlarmZ0Z_5 ;
    wire \Lab_UT.dictrl.nextState_al_1 ;
    wire \Lab_UT.dictrl.nextState_al_1_cascade_ ;
    wire \Lab_UT.dictrl.un2_dicAlarmTrig_i_6 ;
    wire \Lab_UT.dictrl.nextState_al_latmux_1 ;
    wire \Lab_UT.dictrl.nextState_al_latmux_1_cascade_ ;
    wire \Lab_UT.dictrl.nextState_alZ0Z_0 ;
    wire \Lab_UT.dictrl.un2_dicAlarmTrig ;
    wire \Lab_UT.dictrl.N_186 ;
    wire \Lab_UT.dictrl.nextState_al_0_0 ;
    wire \Lab_UT.dictrl.N_186_cascade_ ;
    wire \Lab_UT.dictrl.nextState_al_1_0_0_1 ;
    wire \Lab_UT.dictrl.currState_alZ0Z_0 ;
    wire \Lab_UT.dictrl.currState_alZ0Z_1 ;
    wire \Lab_UT.dictrl.currState_i_5_1 ;
    wire \Lab_UT.dictrl.currState_i_5_0 ;
    wire \Lab_UT.dictrl.un1_currState_8_u_ns_1_cascade_ ;
    wire \Lab_UT.dictrl.currState_ret_7_RNI03VHZ0Z1 ;
    wire \Lab_UT.dictrl.un1_currState_inv_1_cascade_ ;
    wire \Lab_UT.dictrl.currState_0_ret_1_RNIPH7FZ0Z1 ;
    wire \Lab_UT.dictrl.r_dicLdMtens14_1 ;
    wire \Lab_UT.dictrl.r_Sone_init5_1 ;
    wire \Lab_UT.dictrl.currStateZ0Z_3 ;
    wire \Lab_UT.dictrl.un1_currState_inv_1 ;
    wire \Lab_UT.dictrl.N_201_cascade_ ;
    wire \Lab_UT.dictrl.currState_2_RNIOB6H1Z0Z_2 ;
    wire \Lab_UT.dictrl.currStateZ0Z_2 ;
    wire \Lab_UT.dictrl.currState_i_5_3 ;
    wire \Lab_UT.dictrl.r_dicRun_r_1 ;
    wire \Lab_UT.dictrl.r_dicLdMtens15_1i ;
    wire rst;
    wire \Lab_UT.dictrl.r_dicLdMtens15_1 ;
    wire \Lab_UT.dictrl.decoder.de_atSignZ0Z_4_cascade_ ;
    wire \Lab_UT.dictrl.de_atSign ;
    wire \Lab_UT.dictrl.de_littleA_2_cascade_ ;
    wire \Lab_UT.dictrl.de_littleL ;
    wire bu_rx_data_5;
    wire \Lab_UT.dictrl.de_littleL_4 ;
    wire bu_rx_data_6;
    wire \Lab_UT.dictrl.g0_4_2 ;
    wire \Lab_UT.dictrl.de_littleA_2 ;
    wire \Lab_UT.dictrl.decoder.de_littleNZ0Z_1_cascade_ ;
    wire Lab_UT_dictrl_decoder_de_cr_2;
    wire \Lab_UT.n_rdy ;
    wire \resetGen.escKeyZ0Z_3 ;
    wire \buart.Z_rx.sample_g ;
    wire bu_rx_data_7;
    wire bu_rx_data_4;
    wire \Lab_UT.dictrl.decoder.de_atSignZ0Z_5 ;
    wire \Lab_UT.uu0.l_precountZ0Z_0 ;
    wire \uu2.un404_ci_0 ;
    wire \uu2.trig_rd_is_det ;
    wire \uu2.r_addrZ0Z_4 ;
    wire \Lab_UT.di_AMtens_0 ;
    wire \Lab_UT.displayAlarmZ0Z_0 ;
    wire \Lab_UT.di_AStens_0 ;
    wire \Lab_UT.display.N_130 ;
    wire \Lab_UT.display.dOutP_0_iv_i_0_0_cascade_ ;
    wire \Lab_UT.display.dOutP_0_iv_i_1_0 ;
    wire L3_tx_data_0;
    wire \Lab_UT.display.N_153 ;
    wire \Lab_UT.displayAlarmZ1Z_2 ;
    wire \Lab_UT.di_AStens_2 ;
    wire \Lab_UT.display.dOutP_0_iv_i_0_2_cascade_ ;
    wire \Lab_UT.display.dOutP_0_iv_i_1_2 ;
    wire L3_tx_data_2;
    wire \Lab_UT.display.un42_dOutP_1 ;
    wire \Lab_UT.display.cnt_RNI1STE1Z0Z_1 ;
    wire \Lab_UT.display.N_151_cascade_ ;
    wire \Lab_UT.di_AMtens_3 ;
    wire \Lab_UT.display.N_124 ;
    wire rst_g;
    wire \Lab_UT.display.N_106 ;
    wire \Lab_UT.display.N_151 ;
    wire \Lab_UT.di_AMtens_2 ;
    wire \Lab_UT.display.N_115 ;
    wire \Lab_UT.di_AStens_1 ;
    wire \Lab_UT.display.N_108_cascade_ ;
    wire \Lab_UT.di_AMones_1 ;
    wire \Lab_UT.display.dOutP_0_iv_i_0_1 ;
    wire \Lab_UT.display.N_152 ;
    wire \Lab_UT.display.cntZ0Z_1 ;
    wire \Lab_UT.display.N_92 ;
    wire \Lab_UT.display.cntZ0Z_2 ;
    wire \Lab_UT.di_AMtens_1 ;
    wire \Lab_UT.display.cntZ0Z_0 ;
    wire \Lab_UT.display.N_112 ;
    wire \Lab_UT.didp.Sones_subtractor.q_RNO_0Z0Z_3_cascade_ ;
    wire \Lab_UT.didp.Sones_subtractor.q_RNO_0_0_2 ;
    wire \Lab_UT.didp.di_Sones_2 ;
    wire \Lab_UT.didp.di_Sones_3 ;
    wire \Lab_UT.didp.Sones_subtractor.un8_Mtens_ce_cascade_ ;
    wire o_One_Sec_Pulse;
    wire uu0_sec_clkD;
    wire oneSecStrb;
    wire \Lab_UT.ld_enable_dicRun ;
    wire \Lab_UT.didp.N_84_cascade_ ;
    wire \Lab_UT.didp.Sones_subtractor.un8_Mtens_ce ;
    wire \Lab_UT.didp.Stens_subtractor.q_RNI775L5_0Z0Z_3 ;
    wire \Lab_UT.didp.Stens_subtractor.q_RNI775L5_0Z0Z_3_cascade_ ;
    wire \Lab_UT.didp.Stens_subtractor.un1_q_c2 ;
    wire \Lab_UT.didp.Stens_subtractor.q_RNI8PD76Z0Z_1 ;
    wire \Lab_UT.ld_enable_Stens ;
    wire \Lab_UT.didp.Stens_subtractor.q_7_i_1_1 ;
    wire \Lab_UT.didp.Mtens_subtractor.q_RNO_0_3_2_cascade_ ;
    wire \Lab_UT.didp.N_83 ;
    wire \Lab_UT.didp.un3_Mtens_rst_cascade_ ;
    wire \Lab_UT.didp.q_RNI775L5_3 ;
    wire \Lab_UT.didp.Mtens_subtractor.un1_q_axb0_cascade_ ;
    wire \Lab_UT.didp.Mtens_ce ;
    wire \Lab_UT.di_Mtens_2 ;
    wire \Lab_UT.didp.Mtens_ce_cascade_ ;
    wire \Lab_UT.didp.Mtens_subtractor.q_RNO_0_2_3_cascade_ ;
    wire \Lab_UT.didp.di_Mtens_3 ;
    wire \Lab_UT.dicLdMones ;
    wire \Lab_UT.dictrl.r_dicLdMtens14 ;
    wire \Lab_UT.dictrl.de_num0to5_1 ;
    wire \Lab_UT.dicLdMtens_latmux_cascade_ ;
    wire \Lab_UT.didp.di_Stens_2 ;
    wire \Lab_UT.didp.di_Stens_3 ;
    wire \Lab_UT.didp.un6_Mtens_ce ;
    wire \Lab_UT.didp.un3_Mtens_rst ;
    wire \Lab_UT.didp.Mtens_subtractor.q_RNO_2Z0Z_1 ;
    wire \Lab_UT.dicLdMtens ;
    wire \Lab_UT.dicLdMtens_latmux ;
    wire \Lab_UT.didp.Mtens_subtractor.N_147 ;
    wire \Lab_UT.didp.Mtens_subtractor.N_87 ;
    wire \Lab_UT.didp.Mtens_subtractor.N_145 ;
    wire \Lab_UT.didp.Mtens_subtractor.un1_q_c2 ;
    wire \Lab_UT.didp.di_Mtens_1 ;
    wire \Lab_UT.didp.q_RNITOVP_1_cascade_ ;
    wire led_c_1;
    wire \Lab_UT.didp.di_Stens_1 ;
    wire \Lab_UT.didp.q_RNI99F11_1 ;
    wire \Lab_UT.dictrl.r_dicLdMtens15 ;
    wire bu_rx_data_rdy;
    wire \Lab_UT.dictrl.de_num_0 ;
    wire \Lab_UT.dicLdMones_latmux ;
    wire \Lab_UT.displayAlarmZ0Z_6 ;
    wire \Lab_UT.alarm_armed ;
    wire \Lab_UT.displayAlarmZ0Z_4 ;
    wire \Lab_UT.alarm_match ;
    wire \Lab_UT.ld_enable_Sones_cascade_ ;
    wire \Lab_UT.didp.Sones_subtractor.q_RNO_1Z0Z_1 ;
    wire \Lab_UT.didp.Sones_subtractor.q_7_i_1_1_cascade_ ;
    wire \Lab_UT.didp.Sones_subtractor.q_RNI775L5_1_3 ;
    wire \Lab_UT.didp.N_82 ;
    wire \Lab_UT.didp.Sones_subtractor.un1_q_axb0_cascade_ ;
    wire \Lab_UT.didp.Sones_subtractor.N_85 ;
    wire \Lab_UT.didp.di_Sones_1 ;
    wire \Lab_UT.didp.N_81 ;
    wire \Lab_UT.didp.Sones_subtractor.un1_q_c2 ;
    wire \Lab_UT.didp.un4_Mtens_ce ;
    wire \Lab_UT.didp.Mones_subtractor.un1_q_axb_0_cascade_ ;
    wire bu_rx_data_0;
    wire bu_rx_data_3;
    wire bu_rx_data_1;
    wire \Lab_UT.didp.N_84 ;
    wire \Lab_UT.didp.Mones_subtractor.q_0_sqmuxa ;
    wire \Lab_UT.didp.Mones_subtractor.q_RNO_0_2_2_cascade_ ;
    wire bu_rx_data_2;
    wire \Lab_UT.didp.q20_0_i ;
    wire bfn_12_9_0_;
    wire \Lab_UT.didp.Mones_subtractor.un1_q_cry_0_s1 ;
    wire CONSTANT_ONE_NET;
    wire \Lab_UT.didp.di_Mones_2 ;
    wire \Lab_UT.didp.Mones_subtractor.un1_q_cry_1_s1_THRU_CO ;
    wire \Lab_UT.didp.Mones_subtractor.un1_q_cry_1_s1 ;
    wire \Lab_UT.didp.di_Mones_3 ;
    wire \Lab_UT.didp.Mones_subtractor.un1_q_cry_2_s1 ;
    wire \Lab_UT.didp.Mones_subtractor.q_RNO_0_1_3 ;
    wire \Lab_UT.didp.Mones_subtractor.un1_q_cry_0_s1_THRU_CO ;
    wire \Lab_UT.didp.Mones_subtractor.N_80 ;
    wire \Lab_UT.didp.di_Mones_1 ;
    wire \Lab_UT.didp.Mones_subtractor.q_RNO_0Z0Z_1 ;
    wire \Lab_UT.didp.di_MtensZ0Z_0 ;
    wire \Lab_UT.didp.di_Mones_0 ;
    wire \Lab_UT.un1_r_Sone_init5_1_0 ;
    wire \Lab_UT.dictrl.N_258_i ;
    wire \Lab_UT.dicLdSones_latmux ;
    wire \Lab_UT.dicLdSones ;
    wire \Lab_UT.didp.di_Sones_0 ;
    wire \Lab_UT.didp.curr_LEDZ0Z_0 ;
    wire \Lab_UT.didp.di_Stens_0 ;
    wire \Lab_UT.didp.q_RNIRMVP_0 ;
    wire \Lab_UT.didp.q_RNI77F11_0_cascade_ ;
    wire \Lab_UT.didp.curr_LEDZ0Z_1 ;
    wire led_c_0;
    wire \Lab_UT.dictrl.un1_nextState_al24_0 ;
    wire \Lab_UT.alarm_off ;
    wire _gnd_net_;
    wire clk_g;
    wire \Lab_UT.dictrl.nextState_al22 ;

    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .TEST_MODE=1'b0;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .PLLOUT_SELECT="GENCLK";
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FILTER_RANGE=3'b001;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FEEDBACK_PATH="SIMPLE";
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FDA_RELATIVE=4'b0000;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FDA_FEEDBACK=4'b0000;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .ENABLE_ICEGATE=1'b0;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DIVR=4'b0000;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DIVQ=3'b110;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DIVF=7'b0111111;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \latticehx1k_pll_inst.latticehx1k_pll_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(\latticehx1k_pll_inst.clk ),
            .REFERENCECLK(N__10939),
            .RESETB(N__28354),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL());
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_0=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .WRITE_MODE=1;
    defparam \uu2.mem0.ram512X8_inst_physical .READ_MODE=1;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_F=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_E=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_D=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_C=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_B=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_A=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_9=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_8=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_7=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_6=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_5=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_4=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_3=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_2=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_1=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    SB_RAM40_4K \uu2.mem0.ram512X8_inst_physical  (
            .RDATA({dangling_wire_0,\uu2.r_data_wire_7 ,dangling_wire_1,\uu2.r_data_wire_6 ,dangling_wire_2,\uu2.r_data_wire_5 ,dangling_wire_3,\uu2.r_data_wire_4 ,dangling_wire_4,\uu2.r_data_wire_3 ,dangling_wire_5,\uu2.r_data_wire_2 ,dangling_wire_6,\uu2.r_data_wire_1 ,dangling_wire_7,\uu2.r_data_wire_0 }),
            .RADDR({dangling_wire_8,dangling_wire_9,N__13390,N__13363,N__13696,N__22806,N__25114,N__13561,N__13669,N__13636,N__13603}),
            .WADDR({dangling_wire_10,dangling_wire_11,N__12634,N__12700,N__14524,N__14536,N__14551,N__16192,N__14563,N__12685,N__18715}),
            .MASK({dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27}),
            .WDATA({dangling_wire_28,dangling_wire_29,dangling_wire_30,N__18844,dangling_wire_31,N__12574,dangling_wire_32,N__12580,dangling_wire_33,N__12559,dangling_wire_34,N__18817,dangling_wire_35,N__12553,dangling_wire_36,N__12655}),
            .RCLKE(),
            .RCLK(N__29462),
            .RE(N__28355),
            .WCLKE(N__18919),
            .WCLK(N__29461),
            .WE(N__18918));
    IO_PAD led_obuf_1_iopad (
            .OE(N__30236),
            .DIN(N__30235),
            .DOUT(N__30234),
            .PACKAGEPIN(led[1]));
    defparam led_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_1_preio (
            .PADOEN(N__30236),
            .PADOUT(N__30235),
            .PADIN(N__30234),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__27889),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuf_3_iopad (
            .OE(N__30227),
            .DIN(N__30226),
            .DOUT(N__30225),
            .PACKAGEPIN(led[3]));
    defparam led_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_3_preio (
            .PADOEN(N__30227),
            .PADOUT(N__30226),
            .PADIN(N__30225),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__23530),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuf_0_iopad (
            .OE(N__30218),
            .DIN(N__30217),
            .DOUT(N__30216),
            .PACKAGEPIN(led[0]));
    defparam led_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_0_preio (
            .PADOEN(N__30218),
            .PADOUT(N__30217),
            .PADIN(N__30216),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__29596),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD \Z_rcxd.Z_io_iopad  (
            .OE(N__30209),
            .DIN(N__30208),
            .DOUT(N__30207),
            .PACKAGEPIN(from_pc));
    defparam \Z_rcxd.Z_io_preio .PIN_TYPE=6'b000000;
    PRE_IO \Z_rcxd.Z_io_preio  (
            .PADOEN(N__30209),
            .PADOUT(N__30208),
            .PADIN(N__30207),
            .CLOCKENABLE(),
            .DOUT1(GNDG0),
            .OUTPUTENABLE(),
            .DIN0(uart_RXD),
            .DOUT0(GNDG0),
            .INPUTCLK(N__29419),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD clk_in_ibuf_iopad (
            .OE(N__30200),
            .DIN(N__30199),
            .DOUT(N__30198),
            .PACKAGEPIN(clk_in));
    defparam clk_in_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam clk_in_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_in_ibuf_preio (
            .PADOEN(N__30200),
            .PADOUT(N__30199),
            .PADIN(N__30198),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(clk_in_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD to_ir_obuf_iopad (
            .OE(N__30191),
            .DIN(N__30190),
            .DOUT(N__30189),
            .PACKAGEPIN(to_ir));
    defparam to_ir_obuf_preio.NEG_TRIGGER=1'b0;
    defparam to_ir_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO to_ir_obuf_preio (
            .PADOEN(N__30191),
            .PADOUT(N__30190),
            .PADIN(N__30189),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_serial_data_obuf_iopad (
            .OE(N__30182),
            .DIN(N__30181),
            .DOUT(N__30180),
            .PACKAGEPIN(o_serial_data));
    defparam o_serial_data_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_serial_data_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_serial_data_obuf_preio (
            .PADOEN(N__30182),
            .PADOUT(N__30181),
            .PADIN(N__30180),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11923),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD sd_obuf_iopad (
            .OE(N__30173),
            .DIN(N__30172),
            .DOUT(N__30171),
            .PACKAGEPIN(sd));
    defparam sd_obuf_preio.NEG_TRIGGER=1'b0;
    defparam sd_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO sd_obuf_preio (
            .PADOEN(N__30173),
            .PADOUT(N__30172),
            .PADIN(N__30171),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuf_2_iopad (
            .OE(N__30164),
            .DIN(N__30163),
            .DOUT(N__30162),
            .PACKAGEPIN(led[2]));
    defparam led_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_2_preio (
            .PADOEN(N__30164),
            .PADOUT(N__30163),
            .PADIN(N__30162),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__23494),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuf_4_iopad (
            .OE(N__30155),
            .DIN(N__30154),
            .DOUT(N__30153),
            .PACKAGEPIN(led[4]));
    defparam led_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_4_preio (
            .PADOEN(N__30155),
            .PADOUT(N__30154),
            .PADIN(N__30153),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    CascadeMux I__7323 (
            .O(N__30136),
            .I(N__30133));
    InMux I__7322 (
            .O(N__30133),
            .I(N__30130));
    LocalMux I__7321 (
            .O(N__30130),
            .I(\Lab_UT.didp.Mones_subtractor.q_RNO_0_1_3 ));
    InMux I__7320 (
            .O(N__30127),
            .I(N__30124));
    LocalMux I__7319 (
            .O(N__30124),
            .I(\Lab_UT.didp.Mones_subtractor.un1_q_cry_0_s1_THRU_CO ));
    InMux I__7318 (
            .O(N__30121),
            .I(N__30113));
    InMux I__7317 (
            .O(N__30120),
            .I(N__30113));
    InMux I__7316 (
            .O(N__30119),
            .I(N__30108));
    InMux I__7315 (
            .O(N__30118),
            .I(N__30108));
    LocalMux I__7314 (
            .O(N__30113),
            .I(N__30104));
    LocalMux I__7313 (
            .O(N__30108),
            .I(N__30101));
    InMux I__7312 (
            .O(N__30107),
            .I(N__30098));
    Span4Mux_v I__7311 (
            .O(N__30104),
            .I(N__30095));
    Span4Mux_s1_h I__7310 (
            .O(N__30101),
            .I(N__30092));
    LocalMux I__7309 (
            .O(N__30098),
            .I(N__30089));
    Odrv4 I__7308 (
            .O(N__30095),
            .I(\Lab_UT.didp.Mones_subtractor.N_80 ));
    Odrv4 I__7307 (
            .O(N__30092),
            .I(\Lab_UT.didp.Mones_subtractor.N_80 ));
    Odrv12 I__7306 (
            .O(N__30089),
            .I(\Lab_UT.didp.Mones_subtractor.N_80 ));
    InMux I__7305 (
            .O(N__30082),
            .I(N__30078));
    InMux I__7304 (
            .O(N__30081),
            .I(N__30075));
    LocalMux I__7303 (
            .O(N__30078),
            .I(N__30069));
    LocalMux I__7302 (
            .O(N__30075),
            .I(N__30066));
    InMux I__7301 (
            .O(N__30074),
            .I(N__30061));
    InMux I__7300 (
            .O(N__30073),
            .I(N__30061));
    InMux I__7299 (
            .O(N__30072),
            .I(N__30058));
    Span4Mux_h I__7298 (
            .O(N__30069),
            .I(N__30055));
    Odrv4 I__7297 (
            .O(N__30066),
            .I(\Lab_UT.didp.di_Mones_1 ));
    LocalMux I__7296 (
            .O(N__30061),
            .I(\Lab_UT.didp.di_Mones_1 ));
    LocalMux I__7295 (
            .O(N__30058),
            .I(\Lab_UT.didp.di_Mones_1 ));
    Odrv4 I__7294 (
            .O(N__30055),
            .I(\Lab_UT.didp.di_Mones_1 ));
    InMux I__7293 (
            .O(N__30046),
            .I(N__30043));
    LocalMux I__7292 (
            .O(N__30043),
            .I(\Lab_UT.didp.Mones_subtractor.q_RNO_0Z0Z_1 ));
    InMux I__7291 (
            .O(N__30040),
            .I(N__30034));
    InMux I__7290 (
            .O(N__30039),
            .I(N__30031));
    InMux I__7289 (
            .O(N__30038),
            .I(N__30024));
    InMux I__7288 (
            .O(N__30037),
            .I(N__30021));
    LocalMux I__7287 (
            .O(N__30034),
            .I(N__30016));
    LocalMux I__7286 (
            .O(N__30031),
            .I(N__30016));
    InMux I__7285 (
            .O(N__30030),
            .I(N__30013));
    InMux I__7284 (
            .O(N__30029),
            .I(N__30006));
    InMux I__7283 (
            .O(N__30028),
            .I(N__30006));
    InMux I__7282 (
            .O(N__30027),
            .I(N__30006));
    LocalMux I__7281 (
            .O(N__30024),
            .I(N__30003));
    LocalMux I__7280 (
            .O(N__30021),
            .I(\Lab_UT.didp.di_MtensZ0Z_0 ));
    Odrv4 I__7279 (
            .O(N__30016),
            .I(\Lab_UT.didp.di_MtensZ0Z_0 ));
    LocalMux I__7278 (
            .O(N__30013),
            .I(\Lab_UT.didp.di_MtensZ0Z_0 ));
    LocalMux I__7277 (
            .O(N__30006),
            .I(\Lab_UT.didp.di_MtensZ0Z_0 ));
    Odrv12 I__7276 (
            .O(N__30003),
            .I(\Lab_UT.didp.di_MtensZ0Z_0 ));
    InMux I__7275 (
            .O(N__29992),
            .I(N__29989));
    LocalMux I__7274 (
            .O(N__29989),
            .I(N__29982));
    InMux I__7273 (
            .O(N__29988),
            .I(N__29977));
    InMux I__7272 (
            .O(N__29987),
            .I(N__29977));
    InMux I__7271 (
            .O(N__29986),
            .I(N__29972));
    InMux I__7270 (
            .O(N__29985),
            .I(N__29972));
    Span4Mux_h I__7269 (
            .O(N__29982),
            .I(N__29969));
    LocalMux I__7268 (
            .O(N__29977),
            .I(\Lab_UT.didp.di_Mones_0 ));
    LocalMux I__7267 (
            .O(N__29972),
            .I(\Lab_UT.didp.di_Mones_0 ));
    Odrv4 I__7266 (
            .O(N__29969),
            .I(\Lab_UT.didp.di_Mones_0 ));
    CascadeMux I__7265 (
            .O(N__29962),
            .I(N__29953));
    InMux I__7264 (
            .O(N__29961),
            .I(N__29945));
    InMux I__7263 (
            .O(N__29960),
            .I(N__29945));
    InMux I__7262 (
            .O(N__29959),
            .I(N__29940));
    InMux I__7261 (
            .O(N__29958),
            .I(N__29940));
    InMux I__7260 (
            .O(N__29957),
            .I(N__29936));
    InMux I__7259 (
            .O(N__29956),
            .I(N__29929));
    InMux I__7258 (
            .O(N__29953),
            .I(N__29929));
    InMux I__7257 (
            .O(N__29952),
            .I(N__29929));
    InMux I__7256 (
            .O(N__29951),
            .I(N__29924));
    InMux I__7255 (
            .O(N__29950),
            .I(N__29924));
    LocalMux I__7254 (
            .O(N__29945),
            .I(N__29921));
    LocalMux I__7253 (
            .O(N__29940),
            .I(N__29918));
    InMux I__7252 (
            .O(N__29939),
            .I(N__29915));
    LocalMux I__7251 (
            .O(N__29936),
            .I(N__29912));
    LocalMux I__7250 (
            .O(N__29929),
            .I(N__29905));
    LocalMux I__7249 (
            .O(N__29924),
            .I(N__29905));
    Span4Mux_v I__7248 (
            .O(N__29921),
            .I(N__29905));
    Span4Mux_s3_h I__7247 (
            .O(N__29918),
            .I(N__29902));
    LocalMux I__7246 (
            .O(N__29915),
            .I(\Lab_UT.un1_r_Sone_init5_1_0 ));
    Odrv12 I__7245 (
            .O(N__29912),
            .I(\Lab_UT.un1_r_Sone_init5_1_0 ));
    Odrv4 I__7244 (
            .O(N__29905),
            .I(\Lab_UT.un1_r_Sone_init5_1_0 ));
    Odrv4 I__7243 (
            .O(N__29902),
            .I(\Lab_UT.un1_r_Sone_init5_1_0 ));
    InMux I__7242 (
            .O(N__29893),
            .I(N__29888));
    InMux I__7241 (
            .O(N__29892),
            .I(N__29883));
    InMux I__7240 (
            .O(N__29891),
            .I(N__29883));
    LocalMux I__7239 (
            .O(N__29888),
            .I(N__29877));
    LocalMux I__7238 (
            .O(N__29883),
            .I(N__29877));
    InMux I__7237 (
            .O(N__29882),
            .I(N__29874));
    Odrv12 I__7236 (
            .O(N__29877),
            .I(\Lab_UT.dictrl.N_258_i ));
    LocalMux I__7235 (
            .O(N__29874),
            .I(\Lab_UT.dictrl.N_258_i ));
    InMux I__7234 (
            .O(N__29869),
            .I(N__29864));
    InMux I__7233 (
            .O(N__29868),
            .I(N__29859));
    InMux I__7232 (
            .O(N__29867),
            .I(N__29859));
    LocalMux I__7231 (
            .O(N__29864),
            .I(N__29854));
    LocalMux I__7230 (
            .O(N__29859),
            .I(N__29854));
    Span4Mux_v I__7229 (
            .O(N__29854),
            .I(N__29851));
    Span4Mux_h I__7228 (
            .O(N__29851),
            .I(N__29848));
    Odrv4 I__7227 (
            .O(N__29848),
            .I(\Lab_UT.dicLdSones_latmux ));
    CascadeMux I__7226 (
            .O(N__29845),
            .I(N__29840));
    CascadeMux I__7225 (
            .O(N__29844),
            .I(N__29837));
    InMux I__7224 (
            .O(N__29843),
            .I(N__29832));
    InMux I__7223 (
            .O(N__29840),
            .I(N__29832));
    InMux I__7222 (
            .O(N__29837),
            .I(N__29829));
    LocalMux I__7221 (
            .O(N__29832),
            .I(N__29826));
    LocalMux I__7220 (
            .O(N__29829),
            .I(\Lab_UT.dicLdSones ));
    Odrv12 I__7219 (
            .O(N__29826),
            .I(\Lab_UT.dicLdSones ));
    InMux I__7218 (
            .O(N__29821),
            .I(N__29817));
    InMux I__7217 (
            .O(N__29820),
            .I(N__29809));
    LocalMux I__7216 (
            .O(N__29817),
            .I(N__29806));
    InMux I__7215 (
            .O(N__29816),
            .I(N__29799));
    InMux I__7214 (
            .O(N__29815),
            .I(N__29799));
    InMux I__7213 (
            .O(N__29814),
            .I(N__29799));
    InMux I__7212 (
            .O(N__29813),
            .I(N__29794));
    InMux I__7211 (
            .O(N__29812),
            .I(N__29794));
    LocalMux I__7210 (
            .O(N__29809),
            .I(N__29791));
    Odrv4 I__7209 (
            .O(N__29806),
            .I(\Lab_UT.didp.di_Sones_0 ));
    LocalMux I__7208 (
            .O(N__29799),
            .I(\Lab_UT.didp.di_Sones_0 ));
    LocalMux I__7207 (
            .O(N__29794),
            .I(\Lab_UT.didp.di_Sones_0 ));
    Odrv12 I__7206 (
            .O(N__29791),
            .I(\Lab_UT.didp.di_Sones_0 ));
    InMux I__7205 (
            .O(N__29782),
            .I(N__29775));
    InMux I__7204 (
            .O(N__29781),
            .I(N__29768));
    InMux I__7203 (
            .O(N__29780),
            .I(N__29768));
    CascadeMux I__7202 (
            .O(N__29779),
            .I(N__29765));
    CascadeMux I__7201 (
            .O(N__29778),
            .I(N__29762));
    LocalMux I__7200 (
            .O(N__29775),
            .I(N__29758));
    InMux I__7199 (
            .O(N__29774),
            .I(N__29755));
    InMux I__7198 (
            .O(N__29773),
            .I(N__29752));
    LocalMux I__7197 (
            .O(N__29768),
            .I(N__29749));
    InMux I__7196 (
            .O(N__29765),
            .I(N__29744));
    InMux I__7195 (
            .O(N__29762),
            .I(N__29744));
    InMux I__7194 (
            .O(N__29761),
            .I(N__29741));
    Span4Mux_v I__7193 (
            .O(N__29758),
            .I(N__29736));
    LocalMux I__7192 (
            .O(N__29755),
            .I(N__29736));
    LocalMux I__7191 (
            .O(N__29752),
            .I(N__29733));
    Span4Mux_s3_h I__7190 (
            .O(N__29749),
            .I(N__29726));
    LocalMux I__7189 (
            .O(N__29744),
            .I(N__29726));
    LocalMux I__7188 (
            .O(N__29741),
            .I(N__29726));
    Span4Mux_v I__7187 (
            .O(N__29736),
            .I(N__29721));
    Span4Mux_v I__7186 (
            .O(N__29733),
            .I(N__29718));
    Span4Mux_v I__7185 (
            .O(N__29726),
            .I(N__29715));
    InMux I__7184 (
            .O(N__29725),
            .I(N__29710));
    InMux I__7183 (
            .O(N__29724),
            .I(N__29710));
    Odrv4 I__7182 (
            .O(N__29721),
            .I(\Lab_UT.didp.curr_LEDZ0Z_0 ));
    Odrv4 I__7181 (
            .O(N__29718),
            .I(\Lab_UT.didp.curr_LEDZ0Z_0 ));
    Odrv4 I__7180 (
            .O(N__29715),
            .I(\Lab_UT.didp.curr_LEDZ0Z_0 ));
    LocalMux I__7179 (
            .O(N__29710),
            .I(\Lab_UT.didp.curr_LEDZ0Z_0 ));
    InMux I__7178 (
            .O(N__29701),
            .I(N__29696));
    InMux I__7177 (
            .O(N__29700),
            .I(N__29693));
    InMux I__7176 (
            .O(N__29699),
            .I(N__29690));
    LocalMux I__7175 (
            .O(N__29696),
            .I(N__29686));
    LocalMux I__7174 (
            .O(N__29693),
            .I(N__29678));
    LocalMux I__7173 (
            .O(N__29690),
            .I(N__29678));
    InMux I__7172 (
            .O(N__29689),
            .I(N__29675));
    Span4Mux_v I__7171 (
            .O(N__29686),
            .I(N__29672));
    InMux I__7170 (
            .O(N__29685),
            .I(N__29665));
    InMux I__7169 (
            .O(N__29684),
            .I(N__29665));
    InMux I__7168 (
            .O(N__29683),
            .I(N__29665));
    Span4Mux_s3_h I__7167 (
            .O(N__29678),
            .I(N__29660));
    LocalMux I__7166 (
            .O(N__29675),
            .I(N__29660));
    Odrv4 I__7165 (
            .O(N__29672),
            .I(\Lab_UT.didp.di_Stens_0 ));
    LocalMux I__7164 (
            .O(N__29665),
            .I(\Lab_UT.didp.di_Stens_0 ));
    Odrv4 I__7163 (
            .O(N__29660),
            .I(\Lab_UT.didp.di_Stens_0 ));
    InMux I__7162 (
            .O(N__29653),
            .I(N__29650));
    LocalMux I__7161 (
            .O(N__29650),
            .I(\Lab_UT.didp.q_RNIRMVP_0 ));
    CascadeMux I__7160 (
            .O(N__29647),
            .I(\Lab_UT.didp.q_RNI77F11_0_cascade_ ));
    InMux I__7159 (
            .O(N__29644),
            .I(N__29641));
    LocalMux I__7158 (
            .O(N__29641),
            .I(N__29638));
    Span4Mux_v I__7157 (
            .O(N__29638),
            .I(N__29634));
    InMux I__7156 (
            .O(N__29637),
            .I(N__29631));
    IoSpan4Mux I__7155 (
            .O(N__29634),
            .I(N__29624));
    LocalMux I__7154 (
            .O(N__29631),
            .I(N__29624));
    InMux I__7153 (
            .O(N__29630),
            .I(N__29619));
    InMux I__7152 (
            .O(N__29629),
            .I(N__29619));
    Span4Mux_s3_h I__7151 (
            .O(N__29624),
            .I(N__29616));
    LocalMux I__7150 (
            .O(N__29619),
            .I(N__29613));
    Span4Mux_v I__7149 (
            .O(N__29616),
            .I(N__29609));
    Span4Mux_v I__7148 (
            .O(N__29613),
            .I(N__29606));
    InMux I__7147 (
            .O(N__29612),
            .I(N__29603));
    Odrv4 I__7146 (
            .O(N__29609),
            .I(\Lab_UT.didp.curr_LEDZ0Z_1 ));
    Odrv4 I__7145 (
            .O(N__29606),
            .I(\Lab_UT.didp.curr_LEDZ0Z_1 ));
    LocalMux I__7144 (
            .O(N__29603),
            .I(\Lab_UT.didp.curr_LEDZ0Z_1 ));
    IoInMux I__7143 (
            .O(N__29596),
            .I(N__29593));
    LocalMux I__7142 (
            .O(N__29593),
            .I(N__29590));
    Span4Mux_s0_h I__7141 (
            .O(N__29590),
            .I(N__29587));
    Odrv4 I__7140 (
            .O(N__29587),
            .I(led_c_0));
    InMux I__7139 (
            .O(N__29584),
            .I(N__29581));
    LocalMux I__7138 (
            .O(N__29581),
            .I(N__29578));
    Span4Mux_s2_h I__7137 (
            .O(N__29578),
            .I(N__29569));
    InMux I__7136 (
            .O(N__29577),
            .I(N__29562));
    InMux I__7135 (
            .O(N__29576),
            .I(N__29562));
    InMux I__7134 (
            .O(N__29575),
            .I(N__29562));
    InMux I__7133 (
            .O(N__29574),
            .I(N__29555));
    InMux I__7132 (
            .O(N__29573),
            .I(N__29555));
    InMux I__7131 (
            .O(N__29572),
            .I(N__29555));
    Odrv4 I__7130 (
            .O(N__29569),
            .I(\Lab_UT.dictrl.un1_nextState_al24_0 ));
    LocalMux I__7129 (
            .O(N__29562),
            .I(\Lab_UT.dictrl.un1_nextState_al24_0 ));
    LocalMux I__7128 (
            .O(N__29555),
            .I(\Lab_UT.dictrl.un1_nextState_al24_0 ));
    InMux I__7127 (
            .O(N__29548),
            .I(N__29541));
    InMux I__7126 (
            .O(N__29547),
            .I(N__29541));
    InMux I__7125 (
            .O(N__29546),
            .I(N__29536));
    LocalMux I__7124 (
            .O(N__29541),
            .I(N__29533));
    InMux I__7123 (
            .O(N__29540),
            .I(N__29529));
    InMux I__7122 (
            .O(N__29539),
            .I(N__29526));
    LocalMux I__7121 (
            .O(N__29536),
            .I(N__29521));
    Span4Mux_h I__7120 (
            .O(N__29533),
            .I(N__29521));
    InMux I__7119 (
            .O(N__29532),
            .I(N__29518));
    LocalMux I__7118 (
            .O(N__29529),
            .I(N__29513));
    LocalMux I__7117 (
            .O(N__29526),
            .I(N__29513));
    Span4Mux_v I__7116 (
            .O(N__29521),
            .I(N__29509));
    LocalMux I__7115 (
            .O(N__29518),
            .I(N__29506));
    Span4Mux_v I__7114 (
            .O(N__29513),
            .I(N__29503));
    InMux I__7113 (
            .O(N__29512),
            .I(N__29500));
    Odrv4 I__7112 (
            .O(N__29509),
            .I(\Lab_UT.alarm_off ));
    Odrv12 I__7111 (
            .O(N__29506),
            .I(\Lab_UT.alarm_off ));
    Odrv4 I__7110 (
            .O(N__29503),
            .I(\Lab_UT.alarm_off ));
    LocalMux I__7109 (
            .O(N__29500),
            .I(\Lab_UT.alarm_off ));
    CascadeMux I__7108 (
            .O(N__29491),
            .I(N__29487));
    InMux I__7107 (
            .O(N__29490),
            .I(N__29484));
    InMux I__7106 (
            .O(N__29487),
            .I(N__29481));
    LocalMux I__7105 (
            .O(N__29484),
            .I(N__29367));
    LocalMux I__7104 (
            .O(N__29481),
            .I(N__29364));
    ClkMux I__7103 (
            .O(N__29480),
            .I(N__29137));
    ClkMux I__7102 (
            .O(N__29479),
            .I(N__29137));
    ClkMux I__7101 (
            .O(N__29478),
            .I(N__29137));
    ClkMux I__7100 (
            .O(N__29477),
            .I(N__29137));
    ClkMux I__7099 (
            .O(N__29476),
            .I(N__29137));
    ClkMux I__7098 (
            .O(N__29475),
            .I(N__29137));
    ClkMux I__7097 (
            .O(N__29474),
            .I(N__29137));
    ClkMux I__7096 (
            .O(N__29473),
            .I(N__29137));
    ClkMux I__7095 (
            .O(N__29472),
            .I(N__29137));
    ClkMux I__7094 (
            .O(N__29471),
            .I(N__29137));
    ClkMux I__7093 (
            .O(N__29470),
            .I(N__29137));
    ClkMux I__7092 (
            .O(N__29469),
            .I(N__29137));
    ClkMux I__7091 (
            .O(N__29468),
            .I(N__29137));
    ClkMux I__7090 (
            .O(N__29467),
            .I(N__29137));
    ClkMux I__7089 (
            .O(N__29466),
            .I(N__29137));
    ClkMux I__7088 (
            .O(N__29465),
            .I(N__29137));
    ClkMux I__7087 (
            .O(N__29464),
            .I(N__29137));
    ClkMux I__7086 (
            .O(N__29463),
            .I(N__29137));
    ClkMux I__7085 (
            .O(N__29462),
            .I(N__29137));
    ClkMux I__7084 (
            .O(N__29461),
            .I(N__29137));
    ClkMux I__7083 (
            .O(N__29460),
            .I(N__29137));
    ClkMux I__7082 (
            .O(N__29459),
            .I(N__29137));
    ClkMux I__7081 (
            .O(N__29458),
            .I(N__29137));
    ClkMux I__7080 (
            .O(N__29457),
            .I(N__29137));
    ClkMux I__7079 (
            .O(N__29456),
            .I(N__29137));
    ClkMux I__7078 (
            .O(N__29455),
            .I(N__29137));
    ClkMux I__7077 (
            .O(N__29454),
            .I(N__29137));
    ClkMux I__7076 (
            .O(N__29453),
            .I(N__29137));
    ClkMux I__7075 (
            .O(N__29452),
            .I(N__29137));
    ClkMux I__7074 (
            .O(N__29451),
            .I(N__29137));
    ClkMux I__7073 (
            .O(N__29450),
            .I(N__29137));
    ClkMux I__7072 (
            .O(N__29449),
            .I(N__29137));
    ClkMux I__7071 (
            .O(N__29448),
            .I(N__29137));
    ClkMux I__7070 (
            .O(N__29447),
            .I(N__29137));
    ClkMux I__7069 (
            .O(N__29446),
            .I(N__29137));
    ClkMux I__7068 (
            .O(N__29445),
            .I(N__29137));
    ClkMux I__7067 (
            .O(N__29444),
            .I(N__29137));
    ClkMux I__7066 (
            .O(N__29443),
            .I(N__29137));
    ClkMux I__7065 (
            .O(N__29442),
            .I(N__29137));
    ClkMux I__7064 (
            .O(N__29441),
            .I(N__29137));
    ClkMux I__7063 (
            .O(N__29440),
            .I(N__29137));
    ClkMux I__7062 (
            .O(N__29439),
            .I(N__29137));
    ClkMux I__7061 (
            .O(N__29438),
            .I(N__29137));
    ClkMux I__7060 (
            .O(N__29437),
            .I(N__29137));
    ClkMux I__7059 (
            .O(N__29436),
            .I(N__29137));
    ClkMux I__7058 (
            .O(N__29435),
            .I(N__29137));
    ClkMux I__7057 (
            .O(N__29434),
            .I(N__29137));
    ClkMux I__7056 (
            .O(N__29433),
            .I(N__29137));
    ClkMux I__7055 (
            .O(N__29432),
            .I(N__29137));
    ClkMux I__7054 (
            .O(N__29431),
            .I(N__29137));
    ClkMux I__7053 (
            .O(N__29430),
            .I(N__29137));
    ClkMux I__7052 (
            .O(N__29429),
            .I(N__29137));
    ClkMux I__7051 (
            .O(N__29428),
            .I(N__29137));
    ClkMux I__7050 (
            .O(N__29427),
            .I(N__29137));
    ClkMux I__7049 (
            .O(N__29426),
            .I(N__29137));
    ClkMux I__7048 (
            .O(N__29425),
            .I(N__29137));
    ClkMux I__7047 (
            .O(N__29424),
            .I(N__29137));
    ClkMux I__7046 (
            .O(N__29423),
            .I(N__29137));
    ClkMux I__7045 (
            .O(N__29422),
            .I(N__29137));
    ClkMux I__7044 (
            .O(N__29421),
            .I(N__29137));
    ClkMux I__7043 (
            .O(N__29420),
            .I(N__29137));
    ClkMux I__7042 (
            .O(N__29419),
            .I(N__29137));
    ClkMux I__7041 (
            .O(N__29418),
            .I(N__29137));
    ClkMux I__7040 (
            .O(N__29417),
            .I(N__29137));
    ClkMux I__7039 (
            .O(N__29416),
            .I(N__29137));
    ClkMux I__7038 (
            .O(N__29415),
            .I(N__29137));
    ClkMux I__7037 (
            .O(N__29414),
            .I(N__29137));
    ClkMux I__7036 (
            .O(N__29413),
            .I(N__29137));
    ClkMux I__7035 (
            .O(N__29412),
            .I(N__29137));
    ClkMux I__7034 (
            .O(N__29411),
            .I(N__29137));
    ClkMux I__7033 (
            .O(N__29410),
            .I(N__29137));
    ClkMux I__7032 (
            .O(N__29409),
            .I(N__29137));
    ClkMux I__7031 (
            .O(N__29408),
            .I(N__29137));
    ClkMux I__7030 (
            .O(N__29407),
            .I(N__29137));
    ClkMux I__7029 (
            .O(N__29406),
            .I(N__29137));
    ClkMux I__7028 (
            .O(N__29405),
            .I(N__29137));
    ClkMux I__7027 (
            .O(N__29404),
            .I(N__29137));
    ClkMux I__7026 (
            .O(N__29403),
            .I(N__29137));
    ClkMux I__7025 (
            .O(N__29402),
            .I(N__29137));
    ClkMux I__7024 (
            .O(N__29401),
            .I(N__29137));
    ClkMux I__7023 (
            .O(N__29400),
            .I(N__29137));
    ClkMux I__7022 (
            .O(N__29399),
            .I(N__29137));
    ClkMux I__7021 (
            .O(N__29398),
            .I(N__29137));
    ClkMux I__7020 (
            .O(N__29397),
            .I(N__29137));
    ClkMux I__7019 (
            .O(N__29396),
            .I(N__29137));
    ClkMux I__7018 (
            .O(N__29395),
            .I(N__29137));
    ClkMux I__7017 (
            .O(N__29394),
            .I(N__29137));
    ClkMux I__7016 (
            .O(N__29393),
            .I(N__29137));
    ClkMux I__7015 (
            .O(N__29392),
            .I(N__29137));
    ClkMux I__7014 (
            .O(N__29391),
            .I(N__29137));
    ClkMux I__7013 (
            .O(N__29390),
            .I(N__29137));
    ClkMux I__7012 (
            .O(N__29389),
            .I(N__29137));
    ClkMux I__7011 (
            .O(N__29388),
            .I(N__29137));
    ClkMux I__7010 (
            .O(N__29387),
            .I(N__29137));
    ClkMux I__7009 (
            .O(N__29386),
            .I(N__29137));
    ClkMux I__7008 (
            .O(N__29385),
            .I(N__29137));
    ClkMux I__7007 (
            .O(N__29384),
            .I(N__29137));
    ClkMux I__7006 (
            .O(N__29383),
            .I(N__29137));
    ClkMux I__7005 (
            .O(N__29382),
            .I(N__29137));
    ClkMux I__7004 (
            .O(N__29381),
            .I(N__29137));
    ClkMux I__7003 (
            .O(N__29380),
            .I(N__29137));
    ClkMux I__7002 (
            .O(N__29379),
            .I(N__29137));
    ClkMux I__7001 (
            .O(N__29378),
            .I(N__29137));
    ClkMux I__7000 (
            .O(N__29377),
            .I(N__29137));
    ClkMux I__6999 (
            .O(N__29376),
            .I(N__29137));
    ClkMux I__6998 (
            .O(N__29375),
            .I(N__29137));
    ClkMux I__6997 (
            .O(N__29374),
            .I(N__29137));
    ClkMux I__6996 (
            .O(N__29373),
            .I(N__29137));
    ClkMux I__6995 (
            .O(N__29372),
            .I(N__29137));
    ClkMux I__6994 (
            .O(N__29371),
            .I(N__29137));
    ClkMux I__6993 (
            .O(N__29370),
            .I(N__29137));
    Glb2LocalMux I__6992 (
            .O(N__29367),
            .I(N__29137));
    Glb2LocalMux I__6991 (
            .O(N__29364),
            .I(N__29137));
    GlobalMux I__6990 (
            .O(N__29137),
            .I(N__29134));
    gio2CtrlBuf I__6989 (
            .O(N__29134),
            .I(clk_g));
    SRMux I__6988 (
            .O(N__29131),
            .I(N__29127));
    CascadeMux I__6987 (
            .O(N__29130),
            .I(N__29123));
    LocalMux I__6986 (
            .O(N__29127),
            .I(N__29120));
    InMux I__6985 (
            .O(N__29126),
            .I(N__29115));
    InMux I__6984 (
            .O(N__29123),
            .I(N__29115));
    Odrv12 I__6983 (
            .O(N__29120),
            .I(\Lab_UT.dictrl.nextState_al22 ));
    LocalMux I__6982 (
            .O(N__29115),
            .I(\Lab_UT.dictrl.nextState_al22 ));
    CascadeMux I__6981 (
            .O(N__29110),
            .I(\Lab_UT.didp.Mones_subtractor.un1_q_axb_0_cascade_ ));
    InMux I__6980 (
            .O(N__29107),
            .I(N__29099));
    CascadeMux I__6979 (
            .O(N__29106),
            .I(N__29094));
    InMux I__6978 (
            .O(N__29105),
            .I(N__29091));
    InMux I__6977 (
            .O(N__29104),
            .I(N__29086));
    InMux I__6976 (
            .O(N__29103),
            .I(N__29086));
    InMux I__6975 (
            .O(N__29102),
            .I(N__29083));
    LocalMux I__6974 (
            .O(N__29099),
            .I(N__29080));
    InMux I__6973 (
            .O(N__29098),
            .I(N__29077));
    InMux I__6972 (
            .O(N__29097),
            .I(N__29074));
    InMux I__6971 (
            .O(N__29094),
            .I(N__29070));
    LocalMux I__6970 (
            .O(N__29091),
            .I(N__29065));
    LocalMux I__6969 (
            .O(N__29086),
            .I(N__29065));
    LocalMux I__6968 (
            .O(N__29083),
            .I(N__29059));
    Span4Mux_s0_h I__6967 (
            .O(N__29080),
            .I(N__29052));
    LocalMux I__6966 (
            .O(N__29077),
            .I(N__29052));
    LocalMux I__6965 (
            .O(N__29074),
            .I(N__29052));
    InMux I__6964 (
            .O(N__29073),
            .I(N__29049));
    LocalMux I__6963 (
            .O(N__29070),
            .I(N__29042));
    Span4Mux_v I__6962 (
            .O(N__29065),
            .I(N__29042));
    InMux I__6961 (
            .O(N__29064),
            .I(N__29035));
    InMux I__6960 (
            .O(N__29063),
            .I(N__29035));
    InMux I__6959 (
            .O(N__29062),
            .I(N__29035));
    Span4Mux_v I__6958 (
            .O(N__29059),
            .I(N__29030));
    Span4Mux_v I__6957 (
            .O(N__29052),
            .I(N__29030));
    LocalMux I__6956 (
            .O(N__29049),
            .I(N__29027));
    CascadeMux I__6955 (
            .O(N__29048),
            .I(N__29023));
    CascadeMux I__6954 (
            .O(N__29047),
            .I(N__29020));
    Span4Mux_v I__6953 (
            .O(N__29042),
            .I(N__29015));
    LocalMux I__6952 (
            .O(N__29035),
            .I(N__29015));
    Span4Mux_h I__6951 (
            .O(N__29030),
            .I(N__29010));
    Span4Mux_h I__6950 (
            .O(N__29027),
            .I(N__29010));
    InMux I__6949 (
            .O(N__29026),
            .I(N__29003));
    InMux I__6948 (
            .O(N__29023),
            .I(N__29003));
    InMux I__6947 (
            .O(N__29020),
            .I(N__29003));
    Odrv4 I__6946 (
            .O(N__29015),
            .I(bu_rx_data_0));
    Odrv4 I__6945 (
            .O(N__29010),
            .I(bu_rx_data_0));
    LocalMux I__6944 (
            .O(N__29003),
            .I(bu_rx_data_0));
    InMux I__6943 (
            .O(N__28996),
            .I(N__28991));
    CascadeMux I__6942 (
            .O(N__28995),
            .I(N__28988));
    CascadeMux I__6941 (
            .O(N__28994),
            .I(N__28975));
    LocalMux I__6940 (
            .O(N__28991),
            .I(N__28971));
    InMux I__6939 (
            .O(N__28988),
            .I(N__28968));
    InMux I__6938 (
            .O(N__28987),
            .I(N__28965));
    InMux I__6937 (
            .O(N__28986),
            .I(N__28957));
    InMux I__6936 (
            .O(N__28985),
            .I(N__28957));
    InMux I__6935 (
            .O(N__28984),
            .I(N__28957));
    InMux I__6934 (
            .O(N__28983),
            .I(N__28954));
    InMux I__6933 (
            .O(N__28982),
            .I(N__28951));
    InMux I__6932 (
            .O(N__28981),
            .I(N__28948));
    InMux I__6931 (
            .O(N__28980),
            .I(N__28944));
    InMux I__6930 (
            .O(N__28979),
            .I(N__28938));
    InMux I__6929 (
            .O(N__28978),
            .I(N__28938));
    InMux I__6928 (
            .O(N__28975),
            .I(N__28935));
    InMux I__6927 (
            .O(N__28974),
            .I(N__28932));
    Span4Mux_v I__6926 (
            .O(N__28971),
            .I(N__28925));
    LocalMux I__6925 (
            .O(N__28968),
            .I(N__28925));
    LocalMux I__6924 (
            .O(N__28965),
            .I(N__28925));
    CascadeMux I__6923 (
            .O(N__28964),
            .I(N__28921));
    LocalMux I__6922 (
            .O(N__28957),
            .I(N__28916));
    LocalMux I__6921 (
            .O(N__28954),
            .I(N__28916));
    LocalMux I__6920 (
            .O(N__28951),
            .I(N__28913));
    LocalMux I__6919 (
            .O(N__28948),
            .I(N__28910));
    CascadeMux I__6918 (
            .O(N__28947),
            .I(N__28907));
    LocalMux I__6917 (
            .O(N__28944),
            .I(N__28902));
    CascadeMux I__6916 (
            .O(N__28943),
            .I(N__28899));
    LocalMux I__6915 (
            .O(N__28938),
            .I(N__28896));
    LocalMux I__6914 (
            .O(N__28935),
            .I(N__28893));
    LocalMux I__6913 (
            .O(N__28932),
            .I(N__28890));
    Span4Mux_h I__6912 (
            .O(N__28925),
            .I(N__28887));
    InMux I__6911 (
            .O(N__28924),
            .I(N__28884));
    InMux I__6910 (
            .O(N__28921),
            .I(N__28881));
    Span4Mux_v I__6909 (
            .O(N__28916),
            .I(N__28878));
    Span4Mux_v I__6908 (
            .O(N__28913),
            .I(N__28873));
    Span4Mux_h I__6907 (
            .O(N__28910),
            .I(N__28873));
    InMux I__6906 (
            .O(N__28907),
            .I(N__28870));
    InMux I__6905 (
            .O(N__28906),
            .I(N__28867));
    InMux I__6904 (
            .O(N__28905),
            .I(N__28864));
    Span12Mux_v I__6903 (
            .O(N__28902),
            .I(N__28861));
    InMux I__6902 (
            .O(N__28899),
            .I(N__28858));
    Span4Mux_v I__6901 (
            .O(N__28896),
            .I(N__28851));
    Span4Mux_v I__6900 (
            .O(N__28893),
            .I(N__28851));
    Span4Mux_s1_v I__6899 (
            .O(N__28890),
            .I(N__28851));
    Span4Mux_v I__6898 (
            .O(N__28887),
            .I(N__28844));
    LocalMux I__6897 (
            .O(N__28884),
            .I(N__28844));
    LocalMux I__6896 (
            .O(N__28881),
            .I(N__28844));
    Span4Mux_v I__6895 (
            .O(N__28878),
            .I(N__28837));
    Span4Mux_h I__6894 (
            .O(N__28873),
            .I(N__28837));
    LocalMux I__6893 (
            .O(N__28870),
            .I(N__28837));
    LocalMux I__6892 (
            .O(N__28867),
            .I(bu_rx_data_3));
    LocalMux I__6891 (
            .O(N__28864),
            .I(bu_rx_data_3));
    Odrv12 I__6890 (
            .O(N__28861),
            .I(bu_rx_data_3));
    LocalMux I__6889 (
            .O(N__28858),
            .I(bu_rx_data_3));
    Odrv4 I__6888 (
            .O(N__28851),
            .I(bu_rx_data_3));
    Odrv4 I__6887 (
            .O(N__28844),
            .I(bu_rx_data_3));
    Odrv4 I__6886 (
            .O(N__28837),
            .I(bu_rx_data_3));
    CascadeMux I__6885 (
            .O(N__28822),
            .I(N__28813));
    InMux I__6884 (
            .O(N__28821),
            .I(N__28809));
    InMux I__6883 (
            .O(N__28820),
            .I(N__28806));
    InMux I__6882 (
            .O(N__28819),
            .I(N__28803));
    InMux I__6881 (
            .O(N__28818),
            .I(N__28800));
    InMux I__6880 (
            .O(N__28817),
            .I(N__28797));
    InMux I__6879 (
            .O(N__28816),
            .I(N__28792));
    InMux I__6878 (
            .O(N__28813),
            .I(N__28789));
    InMux I__6877 (
            .O(N__28812),
            .I(N__28786));
    LocalMux I__6876 (
            .O(N__28809),
            .I(N__28783));
    LocalMux I__6875 (
            .O(N__28806),
            .I(N__28776));
    LocalMux I__6874 (
            .O(N__28803),
            .I(N__28776));
    LocalMux I__6873 (
            .O(N__28800),
            .I(N__28776));
    LocalMux I__6872 (
            .O(N__28797),
            .I(N__28773));
    InMux I__6871 (
            .O(N__28796),
            .I(N__28766));
    InMux I__6870 (
            .O(N__28795),
            .I(N__28766));
    LocalMux I__6869 (
            .O(N__28792),
            .I(N__28763));
    LocalMux I__6868 (
            .O(N__28789),
            .I(N__28760));
    LocalMux I__6867 (
            .O(N__28786),
            .I(N__28757));
    Span4Mux_v I__6866 (
            .O(N__28783),
            .I(N__28750));
    Span4Mux_v I__6865 (
            .O(N__28776),
            .I(N__28747));
    Span4Mux_s2_v I__6864 (
            .O(N__28773),
            .I(N__28744));
    InMux I__6863 (
            .O(N__28772),
            .I(N__28738));
    InMux I__6862 (
            .O(N__28771),
            .I(N__28738));
    LocalMux I__6861 (
            .O(N__28766),
            .I(N__28735));
    Span4Mux_v I__6860 (
            .O(N__28763),
            .I(N__28732));
    Span4Mux_s2_h I__6859 (
            .O(N__28760),
            .I(N__28729));
    Span12Mux_s8_h I__6858 (
            .O(N__28757),
            .I(N__28726));
    InMux I__6857 (
            .O(N__28756),
            .I(N__28721));
    InMux I__6856 (
            .O(N__28755),
            .I(N__28721));
    InMux I__6855 (
            .O(N__28754),
            .I(N__28718));
    InMux I__6854 (
            .O(N__28753),
            .I(N__28715));
    Span4Mux_v I__6853 (
            .O(N__28750),
            .I(N__28708));
    Span4Mux_v I__6852 (
            .O(N__28747),
            .I(N__28708));
    Span4Mux_h I__6851 (
            .O(N__28744),
            .I(N__28708));
    InMux I__6850 (
            .O(N__28743),
            .I(N__28705));
    LocalMux I__6849 (
            .O(N__28738),
            .I(bu_rx_data_1));
    Odrv12 I__6848 (
            .O(N__28735),
            .I(bu_rx_data_1));
    Odrv4 I__6847 (
            .O(N__28732),
            .I(bu_rx_data_1));
    Odrv4 I__6846 (
            .O(N__28729),
            .I(bu_rx_data_1));
    Odrv12 I__6845 (
            .O(N__28726),
            .I(bu_rx_data_1));
    LocalMux I__6844 (
            .O(N__28721),
            .I(bu_rx_data_1));
    LocalMux I__6843 (
            .O(N__28718),
            .I(bu_rx_data_1));
    LocalMux I__6842 (
            .O(N__28715),
            .I(bu_rx_data_1));
    Odrv4 I__6841 (
            .O(N__28708),
            .I(bu_rx_data_1));
    LocalMux I__6840 (
            .O(N__28705),
            .I(bu_rx_data_1));
    InMux I__6839 (
            .O(N__28684),
            .I(N__28679));
    InMux I__6838 (
            .O(N__28683),
            .I(N__28672));
    InMux I__6837 (
            .O(N__28682),
            .I(N__28672));
    LocalMux I__6836 (
            .O(N__28679),
            .I(N__28669));
    InMux I__6835 (
            .O(N__28678),
            .I(N__28666));
    CascadeMux I__6834 (
            .O(N__28677),
            .I(N__28661));
    LocalMux I__6833 (
            .O(N__28672),
            .I(N__28653));
    Span4Mux_v I__6832 (
            .O(N__28669),
            .I(N__28653));
    LocalMux I__6831 (
            .O(N__28666),
            .I(N__28653));
    InMux I__6830 (
            .O(N__28665),
            .I(N__28644));
    InMux I__6829 (
            .O(N__28664),
            .I(N__28644));
    InMux I__6828 (
            .O(N__28661),
            .I(N__28644));
    InMux I__6827 (
            .O(N__28660),
            .I(N__28644));
    Span4Mux_v I__6826 (
            .O(N__28653),
            .I(N__28641));
    LocalMux I__6825 (
            .O(N__28644),
            .I(\Lab_UT.didp.N_84 ));
    Odrv4 I__6824 (
            .O(N__28641),
            .I(\Lab_UT.didp.N_84 ));
    InMux I__6823 (
            .O(N__28636),
            .I(N__28624));
    InMux I__6822 (
            .O(N__28635),
            .I(N__28624));
    InMux I__6821 (
            .O(N__28634),
            .I(N__28624));
    InMux I__6820 (
            .O(N__28633),
            .I(N__28624));
    LocalMux I__6819 (
            .O(N__28624),
            .I(N__28621));
    Odrv4 I__6818 (
            .O(N__28621),
            .I(\Lab_UT.didp.Mones_subtractor.q_0_sqmuxa ));
    CascadeMux I__6817 (
            .O(N__28618),
            .I(\Lab_UT.didp.Mones_subtractor.q_RNO_0_2_2_cascade_ ));
    InMux I__6816 (
            .O(N__28615),
            .I(N__28603));
    InMux I__6815 (
            .O(N__28614),
            .I(N__28598));
    InMux I__6814 (
            .O(N__28613),
            .I(N__28593));
    CascadeMux I__6813 (
            .O(N__28612),
            .I(N__28590));
    InMux I__6812 (
            .O(N__28611),
            .I(N__28585));
    InMux I__6811 (
            .O(N__28610),
            .I(N__28585));
    InMux I__6810 (
            .O(N__28609),
            .I(N__28580));
    InMux I__6809 (
            .O(N__28608),
            .I(N__28580));
    InMux I__6808 (
            .O(N__28607),
            .I(N__28577));
    InMux I__6807 (
            .O(N__28606),
            .I(N__28574));
    LocalMux I__6806 (
            .O(N__28603),
            .I(N__28570));
    InMux I__6805 (
            .O(N__28602),
            .I(N__28567));
    InMux I__6804 (
            .O(N__28601),
            .I(N__28564));
    LocalMux I__6803 (
            .O(N__28598),
            .I(N__28560));
    InMux I__6802 (
            .O(N__28597),
            .I(N__28557));
    InMux I__6801 (
            .O(N__28596),
            .I(N__28554));
    LocalMux I__6800 (
            .O(N__28593),
            .I(N__28551));
    InMux I__6799 (
            .O(N__28590),
            .I(N__28548));
    LocalMux I__6798 (
            .O(N__28585),
            .I(N__28543));
    LocalMux I__6797 (
            .O(N__28580),
            .I(N__28543));
    LocalMux I__6796 (
            .O(N__28577),
            .I(N__28540));
    LocalMux I__6795 (
            .O(N__28574),
            .I(N__28536));
    InMux I__6794 (
            .O(N__28573),
            .I(N__28533));
    Span4Mux_v I__6793 (
            .O(N__28570),
            .I(N__28530));
    LocalMux I__6792 (
            .O(N__28567),
            .I(N__28527));
    LocalMux I__6791 (
            .O(N__28564),
            .I(N__28524));
    InMux I__6790 (
            .O(N__28563),
            .I(N__28521));
    Span4Mux_v I__6789 (
            .O(N__28560),
            .I(N__28518));
    LocalMux I__6788 (
            .O(N__28557),
            .I(N__28515));
    LocalMux I__6787 (
            .O(N__28554),
            .I(N__28510));
    Span4Mux_s2_v I__6786 (
            .O(N__28551),
            .I(N__28510));
    LocalMux I__6785 (
            .O(N__28548),
            .I(N__28500));
    Span12Mux_s7_v I__6784 (
            .O(N__28543),
            .I(N__28500));
    Span12Mux_s3_h I__6783 (
            .O(N__28540),
            .I(N__28500));
    InMux I__6782 (
            .O(N__28539),
            .I(N__28497));
    Span4Mux_h I__6781 (
            .O(N__28536),
            .I(N__28494));
    LocalMux I__6780 (
            .O(N__28533),
            .I(N__28485));
    Span4Mux_v I__6779 (
            .O(N__28530),
            .I(N__28485));
    Span4Mux_v I__6778 (
            .O(N__28527),
            .I(N__28485));
    Span4Mux_s2_v I__6777 (
            .O(N__28524),
            .I(N__28485));
    LocalMux I__6776 (
            .O(N__28521),
            .I(N__28476));
    Span4Mux_v I__6775 (
            .O(N__28518),
            .I(N__28476));
    Span4Mux_s2_v I__6774 (
            .O(N__28515),
            .I(N__28476));
    Span4Mux_h I__6773 (
            .O(N__28510),
            .I(N__28476));
    InMux I__6772 (
            .O(N__28509),
            .I(N__28469));
    InMux I__6771 (
            .O(N__28508),
            .I(N__28469));
    InMux I__6770 (
            .O(N__28507),
            .I(N__28469));
    Odrv12 I__6769 (
            .O(N__28500),
            .I(bu_rx_data_2));
    LocalMux I__6768 (
            .O(N__28497),
            .I(bu_rx_data_2));
    Odrv4 I__6767 (
            .O(N__28494),
            .I(bu_rx_data_2));
    Odrv4 I__6766 (
            .O(N__28485),
            .I(bu_rx_data_2));
    Odrv4 I__6765 (
            .O(N__28476),
            .I(bu_rx_data_2));
    LocalMux I__6764 (
            .O(N__28469),
            .I(bu_rx_data_2));
    SRMux I__6763 (
            .O(N__28456),
            .I(N__28452));
    SRMux I__6762 (
            .O(N__28455),
            .I(N__28449));
    LocalMux I__6761 (
            .O(N__28452),
            .I(N__28443));
    LocalMux I__6760 (
            .O(N__28449),
            .I(N__28440));
    SRMux I__6759 (
            .O(N__28448),
            .I(N__28437));
    SRMux I__6758 (
            .O(N__28447),
            .I(N__28433));
    SRMux I__6757 (
            .O(N__28446),
            .I(N__28430));
    Span4Mux_s3_h I__6756 (
            .O(N__28443),
            .I(N__28423));
    Span4Mux_s3_h I__6755 (
            .O(N__28440),
            .I(N__28423));
    LocalMux I__6754 (
            .O(N__28437),
            .I(N__28423));
    SRMux I__6753 (
            .O(N__28436),
            .I(N__28420));
    LocalMux I__6752 (
            .O(N__28433),
            .I(N__28416));
    LocalMux I__6751 (
            .O(N__28430),
            .I(N__28413));
    Span4Mux_v I__6750 (
            .O(N__28423),
            .I(N__28408));
    LocalMux I__6749 (
            .O(N__28420),
            .I(N__28408));
    SRMux I__6748 (
            .O(N__28419),
            .I(N__28405));
    Span4Mux_v I__6747 (
            .O(N__28416),
            .I(N__28402));
    Span4Mux_s3_h I__6746 (
            .O(N__28413),
            .I(N__28399));
    Span4Mux_s3_h I__6745 (
            .O(N__28408),
            .I(N__28396));
    LocalMux I__6744 (
            .O(N__28405),
            .I(N__28393));
    Span4Mux_h I__6743 (
            .O(N__28402),
            .I(N__28390));
    Span4Mux_h I__6742 (
            .O(N__28399),
            .I(N__28387));
    Span4Mux_h I__6741 (
            .O(N__28396),
            .I(N__28384));
    Span4Mux_s3_h I__6740 (
            .O(N__28393),
            .I(N__28381));
    Span4Mux_h I__6739 (
            .O(N__28390),
            .I(N__28378));
    Span4Mux_v I__6738 (
            .O(N__28387),
            .I(N__28375));
    Span4Mux_v I__6737 (
            .O(N__28384),
            .I(N__28372));
    Span4Mux_h I__6736 (
            .O(N__28381),
            .I(N__28369));
    Odrv4 I__6735 (
            .O(N__28378),
            .I(\Lab_UT.didp.q20_0_i ));
    Odrv4 I__6734 (
            .O(N__28375),
            .I(\Lab_UT.didp.q20_0_i ));
    Odrv4 I__6733 (
            .O(N__28372),
            .I(\Lab_UT.didp.q20_0_i ));
    Odrv4 I__6732 (
            .O(N__28369),
            .I(\Lab_UT.didp.q20_0_i ));
    InMux I__6731 (
            .O(N__28360),
            .I(\Lab_UT.didp.Mones_subtractor.un1_q_cry_0_s1 ));
    CascadeMux I__6730 (
            .O(N__28357),
            .I(N__28350));
    CascadeMux I__6729 (
            .O(N__28356),
            .I(N__28347));
    SRMux I__6728 (
            .O(N__28355),
            .I(N__28344));
    IoInMux I__6727 (
            .O(N__28354),
            .I(N__28341));
    InMux I__6726 (
            .O(N__28353),
            .I(N__28336));
    InMux I__6725 (
            .O(N__28350),
            .I(N__28336));
    InMux I__6724 (
            .O(N__28347),
            .I(N__28333));
    LocalMux I__6723 (
            .O(N__28344),
            .I(N__28330));
    LocalMux I__6722 (
            .O(N__28341),
            .I(N__28327));
    LocalMux I__6721 (
            .O(N__28336),
            .I(N__28324));
    LocalMux I__6720 (
            .O(N__28333),
            .I(N__28321));
    Span4Mux_h I__6719 (
            .O(N__28330),
            .I(N__28318));
    Span4Mux_s3_v I__6718 (
            .O(N__28327),
            .I(N__28315));
    Span12Mux_s6_h I__6717 (
            .O(N__28324),
            .I(N__28312));
    Span12Mux_s11_v I__6716 (
            .O(N__28321),
            .I(N__28309));
    Span4Mux_h I__6715 (
            .O(N__28318),
            .I(N__28304));
    Span4Mux_h I__6714 (
            .O(N__28315),
            .I(N__28304));
    Odrv12 I__6713 (
            .O(N__28312),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__6712 (
            .O(N__28309),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__6711 (
            .O(N__28304),
            .I(CONSTANT_ONE_NET));
    InMux I__6710 (
            .O(N__28297),
            .I(N__28290));
    InMux I__6709 (
            .O(N__28296),
            .I(N__28290));
    CascadeMux I__6708 (
            .O(N__28295),
            .I(N__28287));
    LocalMux I__6707 (
            .O(N__28290),
            .I(N__28282));
    InMux I__6706 (
            .O(N__28287),
            .I(N__28279));
    InMux I__6705 (
            .O(N__28286),
            .I(N__28274));
    InMux I__6704 (
            .O(N__28285),
            .I(N__28274));
    Sp12to4 I__6703 (
            .O(N__28282),
            .I(N__28271));
    LocalMux I__6702 (
            .O(N__28279),
            .I(\Lab_UT.didp.di_Mones_2 ));
    LocalMux I__6701 (
            .O(N__28274),
            .I(\Lab_UT.didp.di_Mones_2 ));
    Odrv12 I__6700 (
            .O(N__28271),
            .I(\Lab_UT.didp.di_Mones_2 ));
    InMux I__6699 (
            .O(N__28264),
            .I(N__28261));
    LocalMux I__6698 (
            .O(N__28261),
            .I(N__28258));
    Odrv4 I__6697 (
            .O(N__28258),
            .I(\Lab_UT.didp.Mones_subtractor.un1_q_cry_1_s1_THRU_CO ));
    InMux I__6696 (
            .O(N__28255),
            .I(\Lab_UT.didp.Mones_subtractor.un1_q_cry_1_s1 ));
    InMux I__6695 (
            .O(N__28252),
            .I(N__28248));
    InMux I__6694 (
            .O(N__28251),
            .I(N__28244));
    LocalMux I__6693 (
            .O(N__28248),
            .I(N__28241));
    CascadeMux I__6692 (
            .O(N__28247),
            .I(N__28237));
    LocalMux I__6691 (
            .O(N__28244),
            .I(N__28234));
    Span4Mux_h I__6690 (
            .O(N__28241),
            .I(N__28231));
    InMux I__6689 (
            .O(N__28240),
            .I(N__28228));
    InMux I__6688 (
            .O(N__28237),
            .I(N__28225));
    Span4Mux_h I__6687 (
            .O(N__28234),
            .I(N__28222));
    Odrv4 I__6686 (
            .O(N__28231),
            .I(\Lab_UT.didp.di_Mones_3 ));
    LocalMux I__6685 (
            .O(N__28228),
            .I(\Lab_UT.didp.di_Mones_3 ));
    LocalMux I__6684 (
            .O(N__28225),
            .I(\Lab_UT.didp.di_Mones_3 ));
    Odrv4 I__6683 (
            .O(N__28222),
            .I(\Lab_UT.didp.di_Mones_3 ));
    InMux I__6682 (
            .O(N__28213),
            .I(\Lab_UT.didp.Mones_subtractor.un1_q_cry_2_s1 ));
    CascadeMux I__6681 (
            .O(N__28210),
            .I(\Lab_UT.ld_enable_Sones_cascade_ ));
    InMux I__6680 (
            .O(N__28207),
            .I(N__28204));
    LocalMux I__6679 (
            .O(N__28204),
            .I(\Lab_UT.didp.Sones_subtractor.q_RNO_1Z0Z_1 ));
    CascadeMux I__6678 (
            .O(N__28201),
            .I(\Lab_UT.didp.Sones_subtractor.q_7_i_1_1_cascade_ ));
    InMux I__6677 (
            .O(N__28198),
            .I(N__28193));
    InMux I__6676 (
            .O(N__28197),
            .I(N__28188));
    InMux I__6675 (
            .O(N__28196),
            .I(N__28188));
    LocalMux I__6674 (
            .O(N__28193),
            .I(N__28185));
    LocalMux I__6673 (
            .O(N__28188),
            .I(\Lab_UT.didp.Sones_subtractor.q_RNI775L5_1_3 ));
    Odrv4 I__6672 (
            .O(N__28185),
            .I(\Lab_UT.didp.Sones_subtractor.q_RNI775L5_1_3 ));
    InMux I__6671 (
            .O(N__28180),
            .I(N__28176));
    InMux I__6670 (
            .O(N__28179),
            .I(N__28168));
    LocalMux I__6669 (
            .O(N__28176),
            .I(N__28165));
    CascadeMux I__6668 (
            .O(N__28175),
            .I(N__28162));
    InMux I__6667 (
            .O(N__28174),
            .I(N__28156));
    InMux I__6666 (
            .O(N__28173),
            .I(N__28156));
    InMux I__6665 (
            .O(N__28172),
            .I(N__28151));
    InMux I__6664 (
            .O(N__28171),
            .I(N__28151));
    LocalMux I__6663 (
            .O(N__28168),
            .I(N__28148));
    Span4Mux_v I__6662 (
            .O(N__28165),
            .I(N__28145));
    InMux I__6661 (
            .O(N__28162),
            .I(N__28140));
    InMux I__6660 (
            .O(N__28161),
            .I(N__28140));
    LocalMux I__6659 (
            .O(N__28156),
            .I(\Lab_UT.didp.N_82 ));
    LocalMux I__6658 (
            .O(N__28151),
            .I(\Lab_UT.didp.N_82 ));
    Odrv4 I__6657 (
            .O(N__28148),
            .I(\Lab_UT.didp.N_82 ));
    Odrv4 I__6656 (
            .O(N__28145),
            .I(\Lab_UT.didp.N_82 ));
    LocalMux I__6655 (
            .O(N__28140),
            .I(\Lab_UT.didp.N_82 ));
    CascadeMux I__6654 (
            .O(N__28129),
            .I(\Lab_UT.didp.Sones_subtractor.un1_q_axb0_cascade_ ));
    InMux I__6653 (
            .O(N__28126),
            .I(N__28120));
    InMux I__6652 (
            .O(N__28125),
            .I(N__28117));
    InMux I__6651 (
            .O(N__28124),
            .I(N__28112));
    InMux I__6650 (
            .O(N__28123),
            .I(N__28112));
    LocalMux I__6649 (
            .O(N__28120),
            .I(\Lab_UT.didp.Sones_subtractor.N_85 ));
    LocalMux I__6648 (
            .O(N__28117),
            .I(\Lab_UT.didp.Sones_subtractor.N_85 ));
    LocalMux I__6647 (
            .O(N__28112),
            .I(\Lab_UT.didp.Sones_subtractor.N_85 ));
    InMux I__6646 (
            .O(N__28105),
            .I(N__28099));
    InMux I__6645 (
            .O(N__28104),
            .I(N__28096));
    CascadeMux I__6644 (
            .O(N__28103),
            .I(N__28093));
    CascadeMux I__6643 (
            .O(N__28102),
            .I(N__28089));
    LocalMux I__6642 (
            .O(N__28099),
            .I(N__28085));
    LocalMux I__6641 (
            .O(N__28096),
            .I(N__28082));
    InMux I__6640 (
            .O(N__28093),
            .I(N__28077));
    InMux I__6639 (
            .O(N__28092),
            .I(N__28077));
    InMux I__6638 (
            .O(N__28089),
            .I(N__28072));
    InMux I__6637 (
            .O(N__28088),
            .I(N__28072));
    Span4Mux_v I__6636 (
            .O(N__28085),
            .I(N__28067));
    Span4Mux_h I__6635 (
            .O(N__28082),
            .I(N__28067));
    LocalMux I__6634 (
            .O(N__28077),
            .I(\Lab_UT.didp.di_Sones_1 ));
    LocalMux I__6633 (
            .O(N__28072),
            .I(\Lab_UT.didp.di_Sones_1 ));
    Odrv4 I__6632 (
            .O(N__28067),
            .I(\Lab_UT.didp.di_Sones_1 ));
    CascadeMux I__6631 (
            .O(N__28060),
            .I(N__28056));
    CascadeMux I__6630 (
            .O(N__28059),
            .I(N__28052));
    InMux I__6629 (
            .O(N__28056),
            .I(N__28040));
    InMux I__6628 (
            .O(N__28055),
            .I(N__28040));
    InMux I__6627 (
            .O(N__28052),
            .I(N__28040));
    InMux I__6626 (
            .O(N__28051),
            .I(N__28040));
    InMux I__6625 (
            .O(N__28050),
            .I(N__28035));
    InMux I__6624 (
            .O(N__28049),
            .I(N__28035));
    LocalMux I__6623 (
            .O(N__28040),
            .I(\Lab_UT.didp.N_81 ));
    LocalMux I__6622 (
            .O(N__28035),
            .I(\Lab_UT.didp.N_81 ));
    InMux I__6621 (
            .O(N__28030),
            .I(N__28027));
    LocalMux I__6620 (
            .O(N__28027),
            .I(\Lab_UT.didp.Sones_subtractor.un1_q_c2 ));
    InMux I__6619 (
            .O(N__28024),
            .I(N__28016));
    InMux I__6618 (
            .O(N__28023),
            .I(N__28013));
    CascadeMux I__6617 (
            .O(N__28022),
            .I(N__28010));
    CascadeMux I__6616 (
            .O(N__28021),
            .I(N__28007));
    InMux I__6615 (
            .O(N__28020),
            .I(N__28002));
    InMux I__6614 (
            .O(N__28019),
            .I(N__28002));
    LocalMux I__6613 (
            .O(N__28016),
            .I(N__27999));
    LocalMux I__6612 (
            .O(N__28013),
            .I(N__27996));
    InMux I__6611 (
            .O(N__28010),
            .I(N__27991));
    InMux I__6610 (
            .O(N__28007),
            .I(N__27991));
    LocalMux I__6609 (
            .O(N__28002),
            .I(\Lab_UT.didp.un4_Mtens_ce ));
    Odrv4 I__6608 (
            .O(N__27999),
            .I(\Lab_UT.didp.un4_Mtens_ce ));
    Odrv4 I__6607 (
            .O(N__27996),
            .I(\Lab_UT.didp.un4_Mtens_ce ));
    LocalMux I__6606 (
            .O(N__27991),
            .I(\Lab_UT.didp.un4_Mtens_ce ));
    InMux I__6605 (
            .O(N__27982),
            .I(N__27972));
    InMux I__6604 (
            .O(N__27981),
            .I(N__27972));
    InMux I__6603 (
            .O(N__27980),
            .I(N__27972));
    InMux I__6602 (
            .O(N__27979),
            .I(N__27969));
    LocalMux I__6601 (
            .O(N__27972),
            .I(\Lab_UT.didp.Mtens_subtractor.N_87 ));
    LocalMux I__6600 (
            .O(N__27969),
            .I(\Lab_UT.didp.Mtens_subtractor.N_87 ));
    InMux I__6599 (
            .O(N__27964),
            .I(N__27961));
    LocalMux I__6598 (
            .O(N__27961),
            .I(\Lab_UT.didp.Mtens_subtractor.N_145 ));
    InMux I__6597 (
            .O(N__27958),
            .I(N__27955));
    LocalMux I__6596 (
            .O(N__27955),
            .I(N__27952));
    Odrv4 I__6595 (
            .O(N__27952),
            .I(\Lab_UT.didp.Mtens_subtractor.un1_q_c2 ));
    CascadeMux I__6594 (
            .O(N__27949),
            .I(N__27944));
    InMux I__6593 (
            .O(N__27948),
            .I(N__27939));
    CascadeMux I__6592 (
            .O(N__27947),
            .I(N__27935));
    InMux I__6591 (
            .O(N__27944),
            .I(N__27931));
    InMux I__6590 (
            .O(N__27943),
            .I(N__27926));
    InMux I__6589 (
            .O(N__27942),
            .I(N__27926));
    LocalMux I__6588 (
            .O(N__27939),
            .I(N__27923));
    InMux I__6587 (
            .O(N__27938),
            .I(N__27920));
    InMux I__6586 (
            .O(N__27935),
            .I(N__27917));
    InMux I__6585 (
            .O(N__27934),
            .I(N__27914));
    LocalMux I__6584 (
            .O(N__27931),
            .I(N__27911));
    LocalMux I__6583 (
            .O(N__27926),
            .I(N__27908));
    Span4Mux_h I__6582 (
            .O(N__27923),
            .I(N__27905));
    LocalMux I__6581 (
            .O(N__27920),
            .I(\Lab_UT.didp.di_Mtens_1 ));
    LocalMux I__6580 (
            .O(N__27917),
            .I(\Lab_UT.didp.di_Mtens_1 ));
    LocalMux I__6579 (
            .O(N__27914),
            .I(\Lab_UT.didp.di_Mtens_1 ));
    Odrv4 I__6578 (
            .O(N__27911),
            .I(\Lab_UT.didp.di_Mtens_1 ));
    Odrv4 I__6577 (
            .O(N__27908),
            .I(\Lab_UT.didp.di_Mtens_1 ));
    Odrv4 I__6576 (
            .O(N__27905),
            .I(\Lab_UT.didp.di_Mtens_1 ));
    CascadeMux I__6575 (
            .O(N__27892),
            .I(\Lab_UT.didp.q_RNITOVP_1_cascade_ ));
    IoInMux I__6574 (
            .O(N__27889),
            .I(N__27886));
    LocalMux I__6573 (
            .O(N__27886),
            .I(N__27883));
    IoSpan4Mux I__6572 (
            .O(N__27883),
            .I(N__27880));
    Odrv4 I__6571 (
            .O(N__27880),
            .I(led_c_1));
    CascadeMux I__6570 (
            .O(N__27877),
            .I(N__27874));
    InMux I__6569 (
            .O(N__27874),
            .I(N__27864));
    InMux I__6568 (
            .O(N__27873),
            .I(N__27864));
    InMux I__6567 (
            .O(N__27872),
            .I(N__27861));
    InMux I__6566 (
            .O(N__27871),
            .I(N__27858));
    InMux I__6565 (
            .O(N__27870),
            .I(N__27855));
    InMux I__6564 (
            .O(N__27869),
            .I(N__27852));
    LocalMux I__6563 (
            .O(N__27864),
            .I(N__27847));
    LocalMux I__6562 (
            .O(N__27861),
            .I(N__27847));
    LocalMux I__6561 (
            .O(N__27858),
            .I(N__27842));
    LocalMux I__6560 (
            .O(N__27855),
            .I(N__27842));
    LocalMux I__6559 (
            .O(N__27852),
            .I(N__27837));
    Span4Mux_h I__6558 (
            .O(N__27847),
            .I(N__27837));
    Odrv12 I__6557 (
            .O(N__27842),
            .I(\Lab_UT.didp.di_Stens_1 ));
    Odrv4 I__6556 (
            .O(N__27837),
            .I(\Lab_UT.didp.di_Stens_1 ));
    InMux I__6555 (
            .O(N__27832),
            .I(N__27829));
    LocalMux I__6554 (
            .O(N__27829),
            .I(\Lab_UT.didp.q_RNI99F11_1 ));
    InMux I__6553 (
            .O(N__27826),
            .I(N__27823));
    LocalMux I__6552 (
            .O(N__27823),
            .I(N__27820));
    Span4Mux_s3_h I__6551 (
            .O(N__27820),
            .I(N__27817));
    Odrv4 I__6550 (
            .O(N__27817),
            .I(\Lab_UT.dictrl.r_dicLdMtens15 ));
    CascadeMux I__6549 (
            .O(N__27814),
            .I(N__27803));
    InMux I__6548 (
            .O(N__27813),
            .I(N__27799));
    InMux I__6547 (
            .O(N__27812),
            .I(N__27796));
    InMux I__6546 (
            .O(N__27811),
            .I(N__27784));
    CascadeMux I__6545 (
            .O(N__27810),
            .I(N__27778));
    InMux I__6544 (
            .O(N__27809),
            .I(N__27774));
    InMux I__6543 (
            .O(N__27808),
            .I(N__27766));
    InMux I__6542 (
            .O(N__27807),
            .I(N__27766));
    InMux I__6541 (
            .O(N__27806),
            .I(N__27766));
    InMux I__6540 (
            .O(N__27803),
            .I(N__27761));
    InMux I__6539 (
            .O(N__27802),
            .I(N__27761));
    LocalMux I__6538 (
            .O(N__27799),
            .I(N__27756));
    LocalMux I__6537 (
            .O(N__27796),
            .I(N__27756));
    InMux I__6536 (
            .O(N__27795),
            .I(N__27749));
    InMux I__6535 (
            .O(N__27794),
            .I(N__27749));
    InMux I__6534 (
            .O(N__27793),
            .I(N__27749));
    InMux I__6533 (
            .O(N__27792),
            .I(N__27740));
    InMux I__6532 (
            .O(N__27791),
            .I(N__27740));
    InMux I__6531 (
            .O(N__27790),
            .I(N__27735));
    InMux I__6530 (
            .O(N__27789),
            .I(N__27735));
    CascadeMux I__6529 (
            .O(N__27788),
            .I(N__27732));
    InMux I__6528 (
            .O(N__27787),
            .I(N__27726));
    LocalMux I__6527 (
            .O(N__27784),
            .I(N__27722));
    InMux I__6526 (
            .O(N__27783),
            .I(N__27717));
    InMux I__6525 (
            .O(N__27782),
            .I(N__27717));
    InMux I__6524 (
            .O(N__27781),
            .I(N__27713));
    InMux I__6523 (
            .O(N__27778),
            .I(N__27705));
    InMux I__6522 (
            .O(N__27777),
            .I(N__27705));
    LocalMux I__6521 (
            .O(N__27774),
            .I(N__27702));
    InMux I__6520 (
            .O(N__27773),
            .I(N__27697));
    LocalMux I__6519 (
            .O(N__27766),
            .I(N__27692));
    LocalMux I__6518 (
            .O(N__27761),
            .I(N__27692));
    Span4Mux_v I__6517 (
            .O(N__27756),
            .I(N__27687));
    LocalMux I__6516 (
            .O(N__27749),
            .I(N__27687));
    InMux I__6515 (
            .O(N__27748),
            .I(N__27684));
    InMux I__6514 (
            .O(N__27747),
            .I(N__27677));
    InMux I__6513 (
            .O(N__27746),
            .I(N__27677));
    InMux I__6512 (
            .O(N__27745),
            .I(N__27677));
    LocalMux I__6511 (
            .O(N__27740),
            .I(N__27672));
    LocalMux I__6510 (
            .O(N__27735),
            .I(N__27672));
    InMux I__6509 (
            .O(N__27732),
            .I(N__27665));
    InMux I__6508 (
            .O(N__27731),
            .I(N__27665));
    InMux I__6507 (
            .O(N__27730),
            .I(N__27665));
    InMux I__6506 (
            .O(N__27729),
            .I(N__27662));
    LocalMux I__6505 (
            .O(N__27726),
            .I(N__27659));
    InMux I__6504 (
            .O(N__27725),
            .I(N__27656));
    Span4Mux_h I__6503 (
            .O(N__27722),
            .I(N__27651));
    LocalMux I__6502 (
            .O(N__27717),
            .I(N__27651));
    InMux I__6501 (
            .O(N__27716),
            .I(N__27648));
    LocalMux I__6500 (
            .O(N__27713),
            .I(N__27640));
    InMux I__6499 (
            .O(N__27712),
            .I(N__27637));
    InMux I__6498 (
            .O(N__27711),
            .I(N__27632));
    InMux I__6497 (
            .O(N__27710),
            .I(N__27632));
    LocalMux I__6496 (
            .O(N__27705),
            .I(N__27629));
    Span4Mux_h I__6495 (
            .O(N__27702),
            .I(N__27626));
    InMux I__6494 (
            .O(N__27701),
            .I(N__27621));
    InMux I__6493 (
            .O(N__27700),
            .I(N__27621));
    LocalMux I__6492 (
            .O(N__27697),
            .I(N__27612));
    Span4Mux_v I__6491 (
            .O(N__27692),
            .I(N__27612));
    Span4Mux_h I__6490 (
            .O(N__27687),
            .I(N__27612));
    LocalMux I__6489 (
            .O(N__27684),
            .I(N__27612));
    LocalMux I__6488 (
            .O(N__27677),
            .I(N__27605));
    Span4Mux_h I__6487 (
            .O(N__27672),
            .I(N__27605));
    LocalMux I__6486 (
            .O(N__27665),
            .I(N__27605));
    LocalMux I__6485 (
            .O(N__27662),
            .I(N__27594));
    Span4Mux_h I__6484 (
            .O(N__27659),
            .I(N__27594));
    LocalMux I__6483 (
            .O(N__27656),
            .I(N__27594));
    Span4Mux_v I__6482 (
            .O(N__27651),
            .I(N__27594));
    LocalMux I__6481 (
            .O(N__27648),
            .I(N__27594));
    InMux I__6480 (
            .O(N__27647),
            .I(N__27583));
    InMux I__6479 (
            .O(N__27646),
            .I(N__27583));
    InMux I__6478 (
            .O(N__27645),
            .I(N__27583));
    InMux I__6477 (
            .O(N__27644),
            .I(N__27583));
    InMux I__6476 (
            .O(N__27643),
            .I(N__27583));
    Odrv4 I__6475 (
            .O(N__27640),
            .I(bu_rx_data_rdy));
    LocalMux I__6474 (
            .O(N__27637),
            .I(bu_rx_data_rdy));
    LocalMux I__6473 (
            .O(N__27632),
            .I(bu_rx_data_rdy));
    Odrv4 I__6472 (
            .O(N__27629),
            .I(bu_rx_data_rdy));
    Odrv4 I__6471 (
            .O(N__27626),
            .I(bu_rx_data_rdy));
    LocalMux I__6470 (
            .O(N__27621),
            .I(bu_rx_data_rdy));
    Odrv4 I__6469 (
            .O(N__27612),
            .I(bu_rx_data_rdy));
    Odrv4 I__6468 (
            .O(N__27605),
            .I(bu_rx_data_rdy));
    Odrv4 I__6467 (
            .O(N__27594),
            .I(bu_rx_data_rdy));
    LocalMux I__6466 (
            .O(N__27583),
            .I(bu_rx_data_rdy));
    InMux I__6465 (
            .O(N__27562),
            .I(N__27556));
    InMux I__6464 (
            .O(N__27561),
            .I(N__27553));
    InMux I__6463 (
            .O(N__27560),
            .I(N__27546));
    InMux I__6462 (
            .O(N__27559),
            .I(N__27546));
    LocalMux I__6461 (
            .O(N__27556),
            .I(N__27538));
    LocalMux I__6460 (
            .O(N__27553),
            .I(N__27535));
    InMux I__6459 (
            .O(N__27552),
            .I(N__27532));
    InMux I__6458 (
            .O(N__27551),
            .I(N__27529));
    LocalMux I__6457 (
            .O(N__27546),
            .I(N__27526));
    InMux I__6456 (
            .O(N__27545),
            .I(N__27521));
    InMux I__6455 (
            .O(N__27544),
            .I(N__27521));
    InMux I__6454 (
            .O(N__27543),
            .I(N__27518));
    InMux I__6453 (
            .O(N__27542),
            .I(N__27512));
    InMux I__6452 (
            .O(N__27541),
            .I(N__27512));
    Span4Mux_v I__6451 (
            .O(N__27538),
            .I(N__27507));
    Span4Mux_v I__6450 (
            .O(N__27535),
            .I(N__27504));
    LocalMux I__6449 (
            .O(N__27532),
            .I(N__27501));
    LocalMux I__6448 (
            .O(N__27529),
            .I(N__27498));
    Span4Mux_v I__6447 (
            .O(N__27526),
            .I(N__27493));
    LocalMux I__6446 (
            .O(N__27521),
            .I(N__27493));
    LocalMux I__6445 (
            .O(N__27518),
            .I(N__27490));
    InMux I__6444 (
            .O(N__27517),
            .I(N__27487));
    LocalMux I__6443 (
            .O(N__27512),
            .I(N__27484));
    CascadeMux I__6442 (
            .O(N__27511),
            .I(N__27479));
    CascadeMux I__6441 (
            .O(N__27510),
            .I(N__27476));
    Span4Mux_h I__6440 (
            .O(N__27507),
            .I(N__27468));
    Span4Mux_s2_h I__6439 (
            .O(N__27504),
            .I(N__27468));
    Span4Mux_v I__6438 (
            .O(N__27501),
            .I(N__27468));
    Span4Mux_v I__6437 (
            .O(N__27498),
            .I(N__27461));
    Span4Mux_h I__6436 (
            .O(N__27493),
            .I(N__27461));
    Span4Mux_s3_h I__6435 (
            .O(N__27490),
            .I(N__27461));
    LocalMux I__6434 (
            .O(N__27487),
            .I(N__27456));
    Span4Mux_s3_h I__6433 (
            .O(N__27484),
            .I(N__27456));
    InMux I__6432 (
            .O(N__27483),
            .I(N__27445));
    InMux I__6431 (
            .O(N__27482),
            .I(N__27445));
    InMux I__6430 (
            .O(N__27479),
            .I(N__27445));
    InMux I__6429 (
            .O(N__27476),
            .I(N__27445));
    InMux I__6428 (
            .O(N__27475),
            .I(N__27445));
    Odrv4 I__6427 (
            .O(N__27468),
            .I(\Lab_UT.dictrl.de_num_0 ));
    Odrv4 I__6426 (
            .O(N__27461),
            .I(\Lab_UT.dictrl.de_num_0 ));
    Odrv4 I__6425 (
            .O(N__27456),
            .I(\Lab_UT.dictrl.de_num_0 ));
    LocalMux I__6424 (
            .O(N__27445),
            .I(\Lab_UT.dictrl.de_num_0 ));
    InMux I__6423 (
            .O(N__27436),
            .I(N__27430));
    InMux I__6422 (
            .O(N__27435),
            .I(N__27430));
    LocalMux I__6421 (
            .O(N__27430),
            .I(N__27427));
    Odrv4 I__6420 (
            .O(N__27427),
            .I(\Lab_UT.dicLdMones_latmux ));
    InMux I__6419 (
            .O(N__27424),
            .I(N__27421));
    LocalMux I__6418 (
            .O(N__27421),
            .I(N__27418));
    Odrv12 I__6417 (
            .O(N__27418),
            .I(\Lab_UT.displayAlarmZ0Z_6 ));
    InMux I__6416 (
            .O(N__27415),
            .I(N__27408));
    InMux I__6415 (
            .O(N__27414),
            .I(N__27408));
    InMux I__6414 (
            .O(N__27413),
            .I(N__27405));
    LocalMux I__6413 (
            .O(N__27408),
            .I(N__27402));
    LocalMux I__6412 (
            .O(N__27405),
            .I(N__27399));
    Span4Mux_s3_h I__6411 (
            .O(N__27402),
            .I(N__27396));
    Span4Mux_s2_h I__6410 (
            .O(N__27399),
            .I(N__27392));
    Span4Mux_v I__6409 (
            .O(N__27396),
            .I(N__27389));
    CascadeMux I__6408 (
            .O(N__27395),
            .I(N__27385));
    Span4Mux_v I__6407 (
            .O(N__27392),
            .I(N__27382));
    Sp12to4 I__6406 (
            .O(N__27389),
            .I(N__27379));
    InMux I__6405 (
            .O(N__27388),
            .I(N__27374));
    InMux I__6404 (
            .O(N__27385),
            .I(N__27374));
    Odrv4 I__6403 (
            .O(N__27382),
            .I(\Lab_UT.alarm_armed ));
    Odrv12 I__6402 (
            .O(N__27379),
            .I(\Lab_UT.alarm_armed ));
    LocalMux I__6401 (
            .O(N__27374),
            .I(\Lab_UT.alarm_armed ));
    InMux I__6400 (
            .O(N__27367),
            .I(N__27364));
    LocalMux I__6399 (
            .O(N__27364),
            .I(N__27361));
    Span4Mux_v I__6398 (
            .O(N__27361),
            .I(N__27358));
    Odrv4 I__6397 (
            .O(N__27358),
            .I(\Lab_UT.displayAlarmZ0Z_4 ));
    InMux I__6396 (
            .O(N__27355),
            .I(N__27346));
    InMux I__6395 (
            .O(N__27354),
            .I(N__27346));
    InMux I__6394 (
            .O(N__27353),
            .I(N__27346));
    LocalMux I__6393 (
            .O(N__27346),
            .I(N__27342));
    InMux I__6392 (
            .O(N__27345),
            .I(N__27338));
    Span4Mux_h I__6391 (
            .O(N__27342),
            .I(N__27335));
    InMux I__6390 (
            .O(N__27341),
            .I(N__27332));
    LocalMux I__6389 (
            .O(N__27338),
            .I(\Lab_UT.alarm_match ));
    Odrv4 I__6388 (
            .O(N__27335),
            .I(\Lab_UT.alarm_match ));
    LocalMux I__6387 (
            .O(N__27332),
            .I(\Lab_UT.alarm_match ));
    CascadeMux I__6386 (
            .O(N__27325),
            .I(N__27321));
    InMux I__6385 (
            .O(N__27324),
            .I(N__27316));
    InMux I__6384 (
            .O(N__27321),
            .I(N__27316));
    LocalMux I__6383 (
            .O(N__27316),
            .I(\Lab_UT.dicLdMones ));
    InMux I__6382 (
            .O(N__27313),
            .I(N__27310));
    LocalMux I__6381 (
            .O(N__27310),
            .I(N__27307));
    Span4Mux_h I__6380 (
            .O(N__27307),
            .I(N__27304));
    Odrv4 I__6379 (
            .O(N__27304),
            .I(\Lab_UT.dictrl.r_dicLdMtens14 ));
    InMux I__6378 (
            .O(N__27301),
            .I(N__27289));
    InMux I__6377 (
            .O(N__27300),
            .I(N__27286));
    InMux I__6376 (
            .O(N__27299),
            .I(N__27281));
    InMux I__6375 (
            .O(N__27298),
            .I(N__27278));
    InMux I__6374 (
            .O(N__27297),
            .I(N__27271));
    InMux I__6373 (
            .O(N__27296),
            .I(N__27271));
    InMux I__6372 (
            .O(N__27295),
            .I(N__27264));
    InMux I__6371 (
            .O(N__27294),
            .I(N__27264));
    InMux I__6370 (
            .O(N__27293),
            .I(N__27264));
    InMux I__6369 (
            .O(N__27292),
            .I(N__27261));
    LocalMux I__6368 (
            .O(N__27289),
            .I(N__27258));
    LocalMux I__6367 (
            .O(N__27286),
            .I(N__27255));
    InMux I__6366 (
            .O(N__27285),
            .I(N__27250));
    InMux I__6365 (
            .O(N__27284),
            .I(N__27250));
    LocalMux I__6364 (
            .O(N__27281),
            .I(N__27243));
    LocalMux I__6363 (
            .O(N__27278),
            .I(N__27240));
    InMux I__6362 (
            .O(N__27277),
            .I(N__27235));
    InMux I__6361 (
            .O(N__27276),
            .I(N__27235));
    LocalMux I__6360 (
            .O(N__27271),
            .I(N__27232));
    LocalMux I__6359 (
            .O(N__27264),
            .I(N__27227));
    LocalMux I__6358 (
            .O(N__27261),
            .I(N__27227));
    Span4Mux_h I__6357 (
            .O(N__27258),
            .I(N__27220));
    Span4Mux_v I__6356 (
            .O(N__27255),
            .I(N__27220));
    LocalMux I__6355 (
            .O(N__27250),
            .I(N__27220));
    InMux I__6354 (
            .O(N__27249),
            .I(N__27213));
    InMux I__6353 (
            .O(N__27248),
            .I(N__27213));
    InMux I__6352 (
            .O(N__27247),
            .I(N__27213));
    InMux I__6351 (
            .O(N__27246),
            .I(N__27206));
    Span4Mux_h I__6350 (
            .O(N__27243),
            .I(N__27201));
    Span4Mux_s3_h I__6349 (
            .O(N__27240),
            .I(N__27201));
    LocalMux I__6348 (
            .O(N__27235),
            .I(N__27194));
    Span4Mux_s3_h I__6347 (
            .O(N__27232),
            .I(N__27194));
    Span4Mux_h I__6346 (
            .O(N__27227),
            .I(N__27194));
    Span4Mux_h I__6345 (
            .O(N__27220),
            .I(N__27189));
    LocalMux I__6344 (
            .O(N__27213),
            .I(N__27189));
    InMux I__6343 (
            .O(N__27212),
            .I(N__27180));
    InMux I__6342 (
            .O(N__27211),
            .I(N__27180));
    InMux I__6341 (
            .O(N__27210),
            .I(N__27180));
    InMux I__6340 (
            .O(N__27209),
            .I(N__27180));
    LocalMux I__6339 (
            .O(N__27206),
            .I(\Lab_UT.dictrl.de_num0to5_1 ));
    Odrv4 I__6338 (
            .O(N__27201),
            .I(\Lab_UT.dictrl.de_num0to5_1 ));
    Odrv4 I__6337 (
            .O(N__27194),
            .I(\Lab_UT.dictrl.de_num0to5_1 ));
    Odrv4 I__6336 (
            .O(N__27189),
            .I(\Lab_UT.dictrl.de_num0to5_1 ));
    LocalMux I__6335 (
            .O(N__27180),
            .I(\Lab_UT.dictrl.de_num0to5_1 ));
    CascadeMux I__6334 (
            .O(N__27169),
            .I(\Lab_UT.dicLdMtens_latmux_cascade_ ));
    InMux I__6333 (
            .O(N__27166),
            .I(N__27163));
    LocalMux I__6332 (
            .O(N__27163),
            .I(N__27156));
    InMux I__6331 (
            .O(N__27162),
            .I(N__27153));
    InMux I__6330 (
            .O(N__27161),
            .I(N__27148));
    InMux I__6329 (
            .O(N__27160),
            .I(N__27148));
    InMux I__6328 (
            .O(N__27159),
            .I(N__27145));
    Span4Mux_s2_h I__6327 (
            .O(N__27156),
            .I(N__27142));
    LocalMux I__6326 (
            .O(N__27153),
            .I(N__27139));
    LocalMux I__6325 (
            .O(N__27148),
            .I(\Lab_UT.didp.di_Stens_2 ));
    LocalMux I__6324 (
            .O(N__27145),
            .I(\Lab_UT.didp.di_Stens_2 ));
    Odrv4 I__6323 (
            .O(N__27142),
            .I(\Lab_UT.didp.di_Stens_2 ));
    Odrv4 I__6322 (
            .O(N__27139),
            .I(\Lab_UT.didp.di_Stens_2 ));
    CascadeMux I__6321 (
            .O(N__27130),
            .I(N__27127));
    InMux I__6320 (
            .O(N__27127),
            .I(N__27123));
    InMux I__6319 (
            .O(N__27126),
            .I(N__27120));
    LocalMux I__6318 (
            .O(N__27123),
            .I(N__27115));
    LocalMux I__6317 (
            .O(N__27120),
            .I(N__27112));
    InMux I__6316 (
            .O(N__27119),
            .I(N__27109));
    InMux I__6315 (
            .O(N__27118),
            .I(N__27106));
    Span4Mux_s2_h I__6314 (
            .O(N__27115),
            .I(N__27103));
    Span4Mux_h I__6313 (
            .O(N__27112),
            .I(N__27100));
    LocalMux I__6312 (
            .O(N__27109),
            .I(\Lab_UT.didp.di_Stens_3 ));
    LocalMux I__6311 (
            .O(N__27106),
            .I(\Lab_UT.didp.di_Stens_3 ));
    Odrv4 I__6310 (
            .O(N__27103),
            .I(\Lab_UT.didp.di_Stens_3 ));
    Odrv4 I__6309 (
            .O(N__27100),
            .I(\Lab_UT.didp.di_Stens_3 ));
    CascadeMux I__6308 (
            .O(N__27091),
            .I(N__27086));
    CascadeMux I__6307 (
            .O(N__27090),
            .I(N__27082));
    CascadeMux I__6306 (
            .O(N__27089),
            .I(N__27078));
    InMux I__6305 (
            .O(N__27086),
            .I(N__27075));
    InMux I__6304 (
            .O(N__27085),
            .I(N__27068));
    InMux I__6303 (
            .O(N__27082),
            .I(N__27068));
    InMux I__6302 (
            .O(N__27081),
            .I(N__27068));
    InMux I__6301 (
            .O(N__27078),
            .I(N__27065));
    LocalMux I__6300 (
            .O(N__27075),
            .I(N__27062));
    LocalMux I__6299 (
            .O(N__27068),
            .I(N__27059));
    LocalMux I__6298 (
            .O(N__27065),
            .I(\Lab_UT.didp.un6_Mtens_ce ));
    Odrv12 I__6297 (
            .O(N__27062),
            .I(\Lab_UT.didp.un6_Mtens_ce ));
    Odrv4 I__6296 (
            .O(N__27059),
            .I(\Lab_UT.didp.un6_Mtens_ce ));
    InMux I__6295 (
            .O(N__27052),
            .I(N__27047));
    InMux I__6294 (
            .O(N__27051),
            .I(N__27040));
    InMux I__6293 (
            .O(N__27050),
            .I(N__27037));
    LocalMux I__6292 (
            .O(N__27047),
            .I(N__27034));
    InMux I__6291 (
            .O(N__27046),
            .I(N__27025));
    InMux I__6290 (
            .O(N__27045),
            .I(N__27025));
    InMux I__6289 (
            .O(N__27044),
            .I(N__27025));
    InMux I__6288 (
            .O(N__27043),
            .I(N__27025));
    LocalMux I__6287 (
            .O(N__27040),
            .I(\Lab_UT.didp.un3_Mtens_rst ));
    LocalMux I__6286 (
            .O(N__27037),
            .I(\Lab_UT.didp.un3_Mtens_rst ));
    Odrv4 I__6285 (
            .O(N__27034),
            .I(\Lab_UT.didp.un3_Mtens_rst ));
    LocalMux I__6284 (
            .O(N__27025),
            .I(\Lab_UT.didp.un3_Mtens_rst ));
    InMux I__6283 (
            .O(N__27016),
            .I(N__27013));
    LocalMux I__6282 (
            .O(N__27013),
            .I(N__27010));
    Odrv4 I__6281 (
            .O(N__27010),
            .I(\Lab_UT.didp.Mtens_subtractor.q_RNO_2Z0Z_1 ));
    CascadeMux I__6280 (
            .O(N__27007),
            .I(N__27003));
    InMux I__6279 (
            .O(N__27006),
            .I(N__26995));
    InMux I__6278 (
            .O(N__27003),
            .I(N__26995));
    InMux I__6277 (
            .O(N__27002),
            .I(N__26995));
    LocalMux I__6276 (
            .O(N__26995),
            .I(\Lab_UT.dicLdMtens ));
    CascadeMux I__6275 (
            .O(N__26992),
            .I(N__26989));
    InMux I__6274 (
            .O(N__26989),
            .I(N__26983));
    InMux I__6273 (
            .O(N__26988),
            .I(N__26983));
    LocalMux I__6272 (
            .O(N__26983),
            .I(\Lab_UT.dicLdMtens_latmux ));
    InMux I__6271 (
            .O(N__26980),
            .I(N__26977));
    LocalMux I__6270 (
            .O(N__26977),
            .I(\Lab_UT.didp.Mtens_subtractor.N_147 ));
    CascadeMux I__6269 (
            .O(N__26974),
            .I(\Lab_UT.didp.Mtens_subtractor.q_RNO_0_3_2_cascade_ ));
    InMux I__6268 (
            .O(N__26971),
            .I(N__26962));
    InMux I__6267 (
            .O(N__26970),
            .I(N__26962));
    InMux I__6266 (
            .O(N__26969),
            .I(N__26962));
    LocalMux I__6265 (
            .O(N__26962),
            .I(N__26957));
    InMux I__6264 (
            .O(N__26961),
            .I(N__26954));
    CascadeMux I__6263 (
            .O(N__26960),
            .I(N__26951));
    Span4Mux_h I__6262 (
            .O(N__26957),
            .I(N__26947));
    LocalMux I__6261 (
            .O(N__26954),
            .I(N__26944));
    InMux I__6260 (
            .O(N__26951),
            .I(N__26939));
    InMux I__6259 (
            .O(N__26950),
            .I(N__26939));
    Odrv4 I__6258 (
            .O(N__26947),
            .I(\Lab_UT.didp.N_83 ));
    Odrv4 I__6257 (
            .O(N__26944),
            .I(\Lab_UT.didp.N_83 ));
    LocalMux I__6256 (
            .O(N__26939),
            .I(\Lab_UT.didp.N_83 ));
    CascadeMux I__6255 (
            .O(N__26932),
            .I(\Lab_UT.didp.un3_Mtens_rst_cascade_ ));
    InMux I__6254 (
            .O(N__26929),
            .I(N__26926));
    LocalMux I__6253 (
            .O(N__26926),
            .I(N__26923));
    Span4Mux_v I__6252 (
            .O(N__26923),
            .I(N__26920));
    Span4Mux_h I__6251 (
            .O(N__26920),
            .I(N__26915));
    InMux I__6250 (
            .O(N__26919),
            .I(N__26910));
    InMux I__6249 (
            .O(N__26918),
            .I(N__26910));
    Span4Mux_h I__6248 (
            .O(N__26915),
            .I(N__26907));
    LocalMux I__6247 (
            .O(N__26910),
            .I(\Lab_UT.didp.q_RNI775L5_3 ));
    Odrv4 I__6246 (
            .O(N__26907),
            .I(\Lab_UT.didp.q_RNI775L5_3 ));
    CascadeMux I__6245 (
            .O(N__26902),
            .I(\Lab_UT.didp.Mtens_subtractor.un1_q_axb0_cascade_ ));
    CascadeMux I__6244 (
            .O(N__26899),
            .I(N__26896));
    InMux I__6243 (
            .O(N__26896),
            .I(N__26893));
    LocalMux I__6242 (
            .O(N__26893),
            .I(\Lab_UT.didp.Mtens_ce ));
    CascadeMux I__6241 (
            .O(N__26890),
            .I(N__26887));
    InMux I__6240 (
            .O(N__26887),
            .I(N__26883));
    InMux I__6239 (
            .O(N__26886),
            .I(N__26880));
    LocalMux I__6238 (
            .O(N__26883),
            .I(N__26877));
    LocalMux I__6237 (
            .O(N__26880),
            .I(N__26874));
    Span4Mux_v I__6236 (
            .O(N__26877),
            .I(N__26867));
    Span4Mux_v I__6235 (
            .O(N__26874),
            .I(N__26864));
    InMux I__6234 (
            .O(N__26873),
            .I(N__26861));
    InMux I__6233 (
            .O(N__26872),
            .I(N__26854));
    InMux I__6232 (
            .O(N__26871),
            .I(N__26854));
    InMux I__6231 (
            .O(N__26870),
            .I(N__26854));
    Span4Mux_h I__6230 (
            .O(N__26867),
            .I(N__26851));
    Sp12to4 I__6229 (
            .O(N__26864),
            .I(N__26846));
    LocalMux I__6228 (
            .O(N__26861),
            .I(N__26846));
    LocalMux I__6227 (
            .O(N__26854),
            .I(\Lab_UT.di_Mtens_2 ));
    Odrv4 I__6226 (
            .O(N__26851),
            .I(\Lab_UT.di_Mtens_2 ));
    Odrv12 I__6225 (
            .O(N__26846),
            .I(\Lab_UT.di_Mtens_2 ));
    CascadeMux I__6224 (
            .O(N__26839),
            .I(\Lab_UT.didp.Mtens_ce_cascade_ ));
    CascadeMux I__6223 (
            .O(N__26836),
            .I(\Lab_UT.didp.Mtens_subtractor.q_RNO_0_2_3_cascade_ ));
    InMux I__6222 (
            .O(N__26833),
            .I(N__26828));
    InMux I__6221 (
            .O(N__26832),
            .I(N__26825));
    CascadeMux I__6220 (
            .O(N__26831),
            .I(N__26821));
    LocalMux I__6219 (
            .O(N__26828),
            .I(N__26818));
    LocalMux I__6218 (
            .O(N__26825),
            .I(N__26815));
    InMux I__6217 (
            .O(N__26824),
            .I(N__26810));
    InMux I__6216 (
            .O(N__26821),
            .I(N__26810));
    Span4Mux_h I__6215 (
            .O(N__26818),
            .I(N__26807));
    Odrv12 I__6214 (
            .O(N__26815),
            .I(\Lab_UT.didp.di_Mtens_3 ));
    LocalMux I__6213 (
            .O(N__26810),
            .I(\Lab_UT.didp.di_Mtens_3 ));
    Odrv4 I__6212 (
            .O(N__26807),
            .I(\Lab_UT.didp.di_Mtens_3 ));
    InMux I__6211 (
            .O(N__26800),
            .I(N__26797));
    LocalMux I__6210 (
            .O(N__26797),
            .I(N__26791));
    InMux I__6209 (
            .O(N__26796),
            .I(N__26786));
    InMux I__6208 (
            .O(N__26795),
            .I(N__26786));
    InMux I__6207 (
            .O(N__26794),
            .I(N__26781));
    Span4Mux_h I__6206 (
            .O(N__26791),
            .I(N__26778));
    LocalMux I__6205 (
            .O(N__26786),
            .I(N__26775));
    InMux I__6204 (
            .O(N__26785),
            .I(N__26770));
    InMux I__6203 (
            .O(N__26784),
            .I(N__26770));
    LocalMux I__6202 (
            .O(N__26781),
            .I(o_One_Sec_Pulse));
    Odrv4 I__6201 (
            .O(N__26778),
            .I(o_One_Sec_Pulse));
    Odrv12 I__6200 (
            .O(N__26775),
            .I(o_One_Sec_Pulse));
    LocalMux I__6199 (
            .O(N__26770),
            .I(o_One_Sec_Pulse));
    InMux I__6198 (
            .O(N__26761),
            .I(N__26757));
    InMux I__6197 (
            .O(N__26760),
            .I(N__26754));
    LocalMux I__6196 (
            .O(N__26757),
            .I(N__26749));
    LocalMux I__6195 (
            .O(N__26754),
            .I(N__26749));
    Span4Mux_s3_h I__6194 (
            .O(N__26749),
            .I(N__26745));
    InMux I__6193 (
            .O(N__26748),
            .I(N__26742));
    Span4Mux_h I__6192 (
            .O(N__26745),
            .I(N__26739));
    LocalMux I__6191 (
            .O(N__26742),
            .I(uu0_sec_clkD));
    Odrv4 I__6190 (
            .O(N__26739),
            .I(uu0_sec_clkD));
    InMux I__6189 (
            .O(N__26734),
            .I(N__26726));
    InMux I__6188 (
            .O(N__26733),
            .I(N__26719));
    InMux I__6187 (
            .O(N__26732),
            .I(N__26719));
    InMux I__6186 (
            .O(N__26731),
            .I(N__26719));
    InMux I__6185 (
            .O(N__26730),
            .I(N__26714));
    InMux I__6184 (
            .O(N__26729),
            .I(N__26714));
    LocalMux I__6183 (
            .O(N__26726),
            .I(N__26710));
    LocalMux I__6182 (
            .O(N__26719),
            .I(N__26705));
    LocalMux I__6181 (
            .O(N__26714),
            .I(N__26705));
    InMux I__6180 (
            .O(N__26713),
            .I(N__26702));
    Span4Mux_h I__6179 (
            .O(N__26710),
            .I(N__26699));
    Span4Mux_v I__6178 (
            .O(N__26705),
            .I(N__26696));
    LocalMux I__6177 (
            .O(N__26702),
            .I(N__26693));
    Span4Mux_v I__6176 (
            .O(N__26699),
            .I(N__26688));
    Span4Mux_h I__6175 (
            .O(N__26696),
            .I(N__26688));
    Span12Mux_s8_h I__6174 (
            .O(N__26693),
            .I(N__26685));
    Odrv4 I__6173 (
            .O(N__26688),
            .I(oneSecStrb));
    Odrv12 I__6172 (
            .O(N__26685),
            .I(oneSecStrb));
    InMux I__6171 (
            .O(N__26680),
            .I(N__26668));
    InMux I__6170 (
            .O(N__26679),
            .I(N__26668));
    InMux I__6169 (
            .O(N__26678),
            .I(N__26668));
    InMux I__6168 (
            .O(N__26677),
            .I(N__26662));
    InMux I__6167 (
            .O(N__26676),
            .I(N__26662));
    InMux I__6166 (
            .O(N__26675),
            .I(N__26659));
    LocalMux I__6165 (
            .O(N__26668),
            .I(N__26656));
    InMux I__6164 (
            .O(N__26667),
            .I(N__26653));
    LocalMux I__6163 (
            .O(N__26662),
            .I(N__26646));
    LocalMux I__6162 (
            .O(N__26659),
            .I(N__26646));
    Span4Mux_s3_h I__6161 (
            .O(N__26656),
            .I(N__26646));
    LocalMux I__6160 (
            .O(N__26653),
            .I(\Lab_UT.ld_enable_dicRun ));
    Odrv4 I__6159 (
            .O(N__26646),
            .I(\Lab_UT.ld_enable_dicRun ));
    CascadeMux I__6158 (
            .O(N__26641),
            .I(\Lab_UT.didp.N_84_cascade_ ));
    InMux I__6157 (
            .O(N__26638),
            .I(N__26631));
    InMux I__6156 (
            .O(N__26637),
            .I(N__26631));
    InMux I__6155 (
            .O(N__26636),
            .I(N__26628));
    LocalMux I__6154 (
            .O(N__26631),
            .I(\Lab_UT.didp.Sones_subtractor.un8_Mtens_ce ));
    LocalMux I__6153 (
            .O(N__26628),
            .I(\Lab_UT.didp.Sones_subtractor.un8_Mtens_ce ));
    InMux I__6152 (
            .O(N__26623),
            .I(N__26611));
    InMux I__6151 (
            .O(N__26622),
            .I(N__26611));
    InMux I__6150 (
            .O(N__26621),
            .I(N__26611));
    InMux I__6149 (
            .O(N__26620),
            .I(N__26611));
    LocalMux I__6148 (
            .O(N__26611),
            .I(N__26608));
    Odrv4 I__6147 (
            .O(N__26608),
            .I(\Lab_UT.didp.Stens_subtractor.q_RNI775L5_0Z0Z_3 ));
    CascadeMux I__6146 (
            .O(N__26605),
            .I(\Lab_UT.didp.Stens_subtractor.q_RNI775L5_0Z0Z_3_cascade_ ));
    CascadeMux I__6145 (
            .O(N__26602),
            .I(N__26599));
    InMux I__6144 (
            .O(N__26599),
            .I(N__26596));
    LocalMux I__6143 (
            .O(N__26596),
            .I(N__26593));
    Odrv4 I__6142 (
            .O(N__26593),
            .I(\Lab_UT.didp.Stens_subtractor.un1_q_c2 ));
    InMux I__6141 (
            .O(N__26590),
            .I(N__26587));
    LocalMux I__6140 (
            .O(N__26587),
            .I(N__26584));
    Span4Mux_v I__6139 (
            .O(N__26584),
            .I(N__26580));
    InMux I__6138 (
            .O(N__26583),
            .I(N__26577));
    IoSpan4Mux I__6137 (
            .O(N__26580),
            .I(N__26572));
    LocalMux I__6136 (
            .O(N__26577),
            .I(N__26572));
    Odrv4 I__6135 (
            .O(N__26572),
            .I(\Lab_UT.didp.Stens_subtractor.q_RNI8PD76Z0Z_1 ));
    InMux I__6134 (
            .O(N__26569),
            .I(N__26566));
    LocalMux I__6133 (
            .O(N__26566),
            .I(N__26562));
    InMux I__6132 (
            .O(N__26565),
            .I(N__26559));
    Span4Mux_v I__6131 (
            .O(N__26562),
            .I(N__26554));
    LocalMux I__6130 (
            .O(N__26559),
            .I(N__26554));
    Odrv4 I__6129 (
            .O(N__26554),
            .I(\Lab_UT.ld_enable_Stens ));
    InMux I__6128 (
            .O(N__26551),
            .I(N__26548));
    LocalMux I__6127 (
            .O(N__26548),
            .I(N__26545));
    Odrv4 I__6126 (
            .O(N__26545),
            .I(\Lab_UT.didp.Stens_subtractor.q_7_i_1_1 ));
    InMux I__6125 (
            .O(N__26542),
            .I(N__26537));
    InMux I__6124 (
            .O(N__26541),
            .I(N__26532));
    InMux I__6123 (
            .O(N__26540),
            .I(N__26532));
    LocalMux I__6122 (
            .O(N__26537),
            .I(N__26527));
    LocalMux I__6121 (
            .O(N__26532),
            .I(N__26527));
    Span4Mux_h I__6120 (
            .O(N__26527),
            .I(N__26523));
    InMux I__6119 (
            .O(N__26526),
            .I(N__26520));
    Odrv4 I__6118 (
            .O(N__26523),
            .I(\Lab_UT.display.N_152 ));
    LocalMux I__6117 (
            .O(N__26520),
            .I(\Lab_UT.display.N_152 ));
    CascadeMux I__6116 (
            .O(N__26515),
            .I(N__26512));
    InMux I__6115 (
            .O(N__26512),
            .I(N__26504));
    InMux I__6114 (
            .O(N__26511),
            .I(N__26504));
    CascadeMux I__6113 (
            .O(N__26510),
            .I(N__26497));
    InMux I__6112 (
            .O(N__26509),
            .I(N__26492));
    LocalMux I__6111 (
            .O(N__26504),
            .I(N__26487));
    InMux I__6110 (
            .O(N__26503),
            .I(N__26483));
    InMux I__6109 (
            .O(N__26502),
            .I(N__26478));
    InMux I__6108 (
            .O(N__26501),
            .I(N__26478));
    InMux I__6107 (
            .O(N__26500),
            .I(N__26469));
    InMux I__6106 (
            .O(N__26497),
            .I(N__26469));
    InMux I__6105 (
            .O(N__26496),
            .I(N__26469));
    InMux I__6104 (
            .O(N__26495),
            .I(N__26469));
    LocalMux I__6103 (
            .O(N__26492),
            .I(N__26466));
    InMux I__6102 (
            .O(N__26491),
            .I(N__26461));
    InMux I__6101 (
            .O(N__26490),
            .I(N__26461));
    Span4Mux_h I__6100 (
            .O(N__26487),
            .I(N__26458));
    InMux I__6099 (
            .O(N__26486),
            .I(N__26455));
    LocalMux I__6098 (
            .O(N__26483),
            .I(\Lab_UT.display.cntZ0Z_1 ));
    LocalMux I__6097 (
            .O(N__26478),
            .I(\Lab_UT.display.cntZ0Z_1 ));
    LocalMux I__6096 (
            .O(N__26469),
            .I(\Lab_UT.display.cntZ0Z_1 ));
    Odrv4 I__6095 (
            .O(N__26466),
            .I(\Lab_UT.display.cntZ0Z_1 ));
    LocalMux I__6094 (
            .O(N__26461),
            .I(\Lab_UT.display.cntZ0Z_1 ));
    Odrv4 I__6093 (
            .O(N__26458),
            .I(\Lab_UT.display.cntZ0Z_1 ));
    LocalMux I__6092 (
            .O(N__26455),
            .I(\Lab_UT.display.cntZ0Z_1 ));
    InMux I__6091 (
            .O(N__26440),
            .I(N__26434));
    InMux I__6090 (
            .O(N__26439),
            .I(N__26434));
    LocalMux I__6089 (
            .O(N__26434),
            .I(N__26431));
    Odrv4 I__6088 (
            .O(N__26431),
            .I(\Lab_UT.display.N_92 ));
    InMux I__6087 (
            .O(N__26428),
            .I(N__26418));
    InMux I__6086 (
            .O(N__26427),
            .I(N__26418));
    InMux I__6085 (
            .O(N__26426),
            .I(N__26418));
    InMux I__6084 (
            .O(N__26425),
            .I(N__26414));
    LocalMux I__6083 (
            .O(N__26418),
            .I(N__26411));
    CascadeMux I__6082 (
            .O(N__26417),
            .I(N__26403));
    LocalMux I__6081 (
            .O(N__26414),
            .I(N__26398));
    Span4Mux_h I__6080 (
            .O(N__26411),
            .I(N__26395));
    InMux I__6079 (
            .O(N__26410),
            .I(N__26386));
    InMux I__6078 (
            .O(N__26409),
            .I(N__26386));
    InMux I__6077 (
            .O(N__26408),
            .I(N__26386));
    InMux I__6076 (
            .O(N__26407),
            .I(N__26386));
    InMux I__6075 (
            .O(N__26406),
            .I(N__26383));
    InMux I__6074 (
            .O(N__26403),
            .I(N__26376));
    InMux I__6073 (
            .O(N__26402),
            .I(N__26376));
    InMux I__6072 (
            .O(N__26401),
            .I(N__26376));
    Odrv4 I__6071 (
            .O(N__26398),
            .I(\Lab_UT.display.cntZ0Z_2 ));
    Odrv4 I__6070 (
            .O(N__26395),
            .I(\Lab_UT.display.cntZ0Z_2 ));
    LocalMux I__6069 (
            .O(N__26386),
            .I(\Lab_UT.display.cntZ0Z_2 ));
    LocalMux I__6068 (
            .O(N__26383),
            .I(\Lab_UT.display.cntZ0Z_2 ));
    LocalMux I__6067 (
            .O(N__26376),
            .I(\Lab_UT.display.cntZ0Z_2 ));
    CascadeMux I__6066 (
            .O(N__26365),
            .I(N__26362));
    InMux I__6065 (
            .O(N__26362),
            .I(N__26359));
    LocalMux I__6064 (
            .O(N__26359),
            .I(N__26356));
    Span4Mux_v I__6063 (
            .O(N__26356),
            .I(N__26351));
    InMux I__6062 (
            .O(N__26355),
            .I(N__26346));
    InMux I__6061 (
            .O(N__26354),
            .I(N__26346));
    Odrv4 I__6060 (
            .O(N__26351),
            .I(\Lab_UT.di_AMtens_1 ));
    LocalMux I__6059 (
            .O(N__26346),
            .I(\Lab_UT.di_AMtens_1 ));
    CascadeMux I__6058 (
            .O(N__26341),
            .I(N__26338));
    InMux I__6057 (
            .O(N__26338),
            .I(N__26328));
    InMux I__6056 (
            .O(N__26337),
            .I(N__26321));
    InMux I__6055 (
            .O(N__26336),
            .I(N__26321));
    InMux I__6054 (
            .O(N__26335),
            .I(N__26321));
    CascadeMux I__6053 (
            .O(N__26334),
            .I(N__26318));
    InMux I__6052 (
            .O(N__26333),
            .I(N__26310));
    InMux I__6051 (
            .O(N__26332),
            .I(N__26310));
    InMux I__6050 (
            .O(N__26331),
            .I(N__26310));
    LocalMux I__6049 (
            .O(N__26328),
            .I(N__26305));
    LocalMux I__6048 (
            .O(N__26321),
            .I(N__26305));
    InMux I__6047 (
            .O(N__26318),
            .I(N__26302));
    CascadeMux I__6046 (
            .O(N__26317),
            .I(N__26294));
    LocalMux I__6045 (
            .O(N__26310),
            .I(N__26289));
    Span4Mux_h I__6044 (
            .O(N__26305),
            .I(N__26284));
    LocalMux I__6043 (
            .O(N__26302),
            .I(N__26284));
    InMux I__6042 (
            .O(N__26301),
            .I(N__26273));
    InMux I__6041 (
            .O(N__26300),
            .I(N__26273));
    InMux I__6040 (
            .O(N__26299),
            .I(N__26273));
    InMux I__6039 (
            .O(N__26298),
            .I(N__26273));
    InMux I__6038 (
            .O(N__26297),
            .I(N__26273));
    InMux I__6037 (
            .O(N__26294),
            .I(N__26266));
    InMux I__6036 (
            .O(N__26293),
            .I(N__26266));
    InMux I__6035 (
            .O(N__26292),
            .I(N__26266));
    Odrv4 I__6034 (
            .O(N__26289),
            .I(\Lab_UT.display.cntZ0Z_0 ));
    Odrv4 I__6033 (
            .O(N__26284),
            .I(\Lab_UT.display.cntZ0Z_0 ));
    LocalMux I__6032 (
            .O(N__26273),
            .I(\Lab_UT.display.cntZ0Z_0 ));
    LocalMux I__6031 (
            .O(N__26266),
            .I(\Lab_UT.display.cntZ0Z_0 ));
    InMux I__6030 (
            .O(N__26257),
            .I(N__26254));
    LocalMux I__6029 (
            .O(N__26254),
            .I(N__26251));
    Span4Mux_h I__6028 (
            .O(N__26251),
            .I(N__26248));
    Odrv4 I__6027 (
            .O(N__26248),
            .I(\Lab_UT.display.N_112 ));
    CascadeMux I__6026 (
            .O(N__26245),
            .I(\Lab_UT.didp.Sones_subtractor.q_RNO_0Z0Z_3_cascade_ ));
    CascadeMux I__6025 (
            .O(N__26242),
            .I(N__26239));
    InMux I__6024 (
            .O(N__26239),
            .I(N__26236));
    LocalMux I__6023 (
            .O(N__26236),
            .I(\Lab_UT.didp.Sones_subtractor.q_RNO_0_0_2 ));
    InMux I__6022 (
            .O(N__26233),
            .I(N__26230));
    LocalMux I__6021 (
            .O(N__26230),
            .I(N__26226));
    InMux I__6020 (
            .O(N__26229),
            .I(N__26220));
    Span4Mux_v I__6019 (
            .O(N__26226),
            .I(N__26217));
    InMux I__6018 (
            .O(N__26225),
            .I(N__26214));
    InMux I__6017 (
            .O(N__26224),
            .I(N__26209));
    InMux I__6016 (
            .O(N__26223),
            .I(N__26209));
    LocalMux I__6015 (
            .O(N__26220),
            .I(N__26206));
    Odrv4 I__6014 (
            .O(N__26217),
            .I(\Lab_UT.didp.di_Sones_2 ));
    LocalMux I__6013 (
            .O(N__26214),
            .I(\Lab_UT.didp.di_Sones_2 ));
    LocalMux I__6012 (
            .O(N__26209),
            .I(\Lab_UT.didp.di_Sones_2 ));
    Odrv4 I__6011 (
            .O(N__26206),
            .I(\Lab_UT.didp.di_Sones_2 ));
    InMux I__6010 (
            .O(N__26197),
            .I(N__26194));
    LocalMux I__6009 (
            .O(N__26194),
            .I(N__26189));
    CascadeMux I__6008 (
            .O(N__26193),
            .I(N__26185));
    CascadeMux I__6007 (
            .O(N__26192),
            .I(N__26182));
    Span4Mux_v I__6006 (
            .O(N__26189),
            .I(N__26179));
    InMux I__6005 (
            .O(N__26188),
            .I(N__26176));
    InMux I__6004 (
            .O(N__26185),
            .I(N__26171));
    InMux I__6003 (
            .O(N__26182),
            .I(N__26171));
    Sp12to4 I__6002 (
            .O(N__26179),
            .I(N__26166));
    LocalMux I__6001 (
            .O(N__26176),
            .I(N__26166));
    LocalMux I__6000 (
            .O(N__26171),
            .I(\Lab_UT.didp.di_Sones_3 ));
    Odrv12 I__5999 (
            .O(N__26166),
            .I(\Lab_UT.didp.di_Sones_3 ));
    CascadeMux I__5998 (
            .O(N__26161),
            .I(\Lab_UT.didp.Sones_subtractor.un8_Mtens_ce_cascade_ ));
    CascadeMux I__5997 (
            .O(N__26158),
            .I(N__26153));
    InMux I__5996 (
            .O(N__26157),
            .I(N__26138));
    InMux I__5995 (
            .O(N__26156),
            .I(N__26138));
    InMux I__5994 (
            .O(N__26153),
            .I(N__26135));
    InMux I__5993 (
            .O(N__26152),
            .I(N__26130));
    InMux I__5992 (
            .O(N__26151),
            .I(N__26130));
    InMux I__5991 (
            .O(N__26150),
            .I(N__26127));
    InMux I__5990 (
            .O(N__26149),
            .I(N__26124));
    InMux I__5989 (
            .O(N__26148),
            .I(N__26121));
    InMux I__5988 (
            .O(N__26147),
            .I(N__26118));
    InMux I__5987 (
            .O(N__26146),
            .I(N__26115));
    InMux I__5986 (
            .O(N__26145),
            .I(N__26110));
    InMux I__5985 (
            .O(N__26144),
            .I(N__26110));
    InMux I__5984 (
            .O(N__26143),
            .I(N__26107));
    LocalMux I__5983 (
            .O(N__26138),
            .I(N__26060));
    LocalMux I__5982 (
            .O(N__26135),
            .I(N__26057));
    LocalMux I__5981 (
            .O(N__26130),
            .I(N__26054));
    LocalMux I__5980 (
            .O(N__26127),
            .I(N__26051));
    LocalMux I__5979 (
            .O(N__26124),
            .I(N__26034));
    LocalMux I__5978 (
            .O(N__26121),
            .I(N__26031));
    LocalMux I__5977 (
            .O(N__26118),
            .I(N__26028));
    LocalMux I__5976 (
            .O(N__26115),
            .I(N__26025));
    LocalMux I__5975 (
            .O(N__26110),
            .I(N__26022));
    LocalMux I__5974 (
            .O(N__26107),
            .I(N__26019));
    SRMux I__5973 (
            .O(N__26106),
            .I(N__25882));
    SRMux I__5972 (
            .O(N__26105),
            .I(N__25882));
    SRMux I__5971 (
            .O(N__26104),
            .I(N__25882));
    SRMux I__5970 (
            .O(N__26103),
            .I(N__25882));
    SRMux I__5969 (
            .O(N__26102),
            .I(N__25882));
    SRMux I__5968 (
            .O(N__26101),
            .I(N__25882));
    SRMux I__5967 (
            .O(N__26100),
            .I(N__25882));
    SRMux I__5966 (
            .O(N__26099),
            .I(N__25882));
    SRMux I__5965 (
            .O(N__26098),
            .I(N__25882));
    SRMux I__5964 (
            .O(N__26097),
            .I(N__25882));
    SRMux I__5963 (
            .O(N__26096),
            .I(N__25882));
    SRMux I__5962 (
            .O(N__26095),
            .I(N__25882));
    SRMux I__5961 (
            .O(N__26094),
            .I(N__25882));
    SRMux I__5960 (
            .O(N__26093),
            .I(N__25882));
    SRMux I__5959 (
            .O(N__26092),
            .I(N__25882));
    SRMux I__5958 (
            .O(N__26091),
            .I(N__25882));
    SRMux I__5957 (
            .O(N__26090),
            .I(N__25882));
    SRMux I__5956 (
            .O(N__26089),
            .I(N__25882));
    SRMux I__5955 (
            .O(N__26088),
            .I(N__25882));
    SRMux I__5954 (
            .O(N__26087),
            .I(N__25882));
    SRMux I__5953 (
            .O(N__26086),
            .I(N__25882));
    SRMux I__5952 (
            .O(N__26085),
            .I(N__25882));
    SRMux I__5951 (
            .O(N__26084),
            .I(N__25882));
    SRMux I__5950 (
            .O(N__26083),
            .I(N__25882));
    SRMux I__5949 (
            .O(N__26082),
            .I(N__25882));
    SRMux I__5948 (
            .O(N__26081),
            .I(N__25882));
    SRMux I__5947 (
            .O(N__26080),
            .I(N__25882));
    SRMux I__5946 (
            .O(N__26079),
            .I(N__25882));
    SRMux I__5945 (
            .O(N__26078),
            .I(N__25882));
    SRMux I__5944 (
            .O(N__26077),
            .I(N__25882));
    SRMux I__5943 (
            .O(N__26076),
            .I(N__25882));
    SRMux I__5942 (
            .O(N__26075),
            .I(N__25882));
    SRMux I__5941 (
            .O(N__26074),
            .I(N__25882));
    SRMux I__5940 (
            .O(N__26073),
            .I(N__25882));
    SRMux I__5939 (
            .O(N__26072),
            .I(N__25882));
    SRMux I__5938 (
            .O(N__26071),
            .I(N__25882));
    SRMux I__5937 (
            .O(N__26070),
            .I(N__25882));
    SRMux I__5936 (
            .O(N__26069),
            .I(N__25882));
    SRMux I__5935 (
            .O(N__26068),
            .I(N__25882));
    SRMux I__5934 (
            .O(N__26067),
            .I(N__25882));
    SRMux I__5933 (
            .O(N__26066),
            .I(N__25882));
    SRMux I__5932 (
            .O(N__26065),
            .I(N__25882));
    SRMux I__5931 (
            .O(N__26064),
            .I(N__25882));
    SRMux I__5930 (
            .O(N__26063),
            .I(N__25882));
    Glb2LocalMux I__5929 (
            .O(N__26060),
            .I(N__25882));
    Glb2LocalMux I__5928 (
            .O(N__26057),
            .I(N__25882));
    Glb2LocalMux I__5927 (
            .O(N__26054),
            .I(N__25882));
    Glb2LocalMux I__5926 (
            .O(N__26051),
            .I(N__25882));
    SRMux I__5925 (
            .O(N__26050),
            .I(N__25882));
    SRMux I__5924 (
            .O(N__26049),
            .I(N__25882));
    SRMux I__5923 (
            .O(N__26048),
            .I(N__25882));
    SRMux I__5922 (
            .O(N__26047),
            .I(N__25882));
    SRMux I__5921 (
            .O(N__26046),
            .I(N__25882));
    SRMux I__5920 (
            .O(N__26045),
            .I(N__25882));
    SRMux I__5919 (
            .O(N__26044),
            .I(N__25882));
    SRMux I__5918 (
            .O(N__26043),
            .I(N__25882));
    SRMux I__5917 (
            .O(N__26042),
            .I(N__25882));
    SRMux I__5916 (
            .O(N__26041),
            .I(N__25882));
    SRMux I__5915 (
            .O(N__26040),
            .I(N__25882));
    SRMux I__5914 (
            .O(N__26039),
            .I(N__25882));
    SRMux I__5913 (
            .O(N__26038),
            .I(N__25882));
    SRMux I__5912 (
            .O(N__26037),
            .I(N__25882));
    Glb2LocalMux I__5911 (
            .O(N__26034),
            .I(N__25882));
    Glb2LocalMux I__5910 (
            .O(N__26031),
            .I(N__25882));
    Glb2LocalMux I__5909 (
            .O(N__26028),
            .I(N__25882));
    Glb2LocalMux I__5908 (
            .O(N__26025),
            .I(N__25882));
    Glb2LocalMux I__5907 (
            .O(N__26022),
            .I(N__25882));
    Glb2LocalMux I__5906 (
            .O(N__26019),
            .I(N__25882));
    GlobalMux I__5905 (
            .O(N__25882),
            .I(N__25879));
    gio2CtrlBuf I__5904 (
            .O(N__25879),
            .I(rst_g));
    InMux I__5903 (
            .O(N__25876),
            .I(N__25870));
    InMux I__5902 (
            .O(N__25875),
            .I(N__25870));
    LocalMux I__5901 (
            .O(N__25870),
            .I(\Lab_UT.display.N_106 ));
    InMux I__5900 (
            .O(N__25867),
            .I(N__25862));
    InMux I__5899 (
            .O(N__25866),
            .I(N__25857));
    InMux I__5898 (
            .O(N__25865),
            .I(N__25857));
    LocalMux I__5897 (
            .O(N__25862),
            .I(\Lab_UT.display.N_151 ));
    LocalMux I__5896 (
            .O(N__25857),
            .I(\Lab_UT.display.N_151 ));
    InMux I__5895 (
            .O(N__25852),
            .I(N__25848));
    InMux I__5894 (
            .O(N__25851),
            .I(N__25845));
    LocalMux I__5893 (
            .O(N__25848),
            .I(N__25840));
    LocalMux I__5892 (
            .O(N__25845),
            .I(N__25837));
    InMux I__5891 (
            .O(N__25844),
            .I(N__25834));
    InMux I__5890 (
            .O(N__25843),
            .I(N__25831));
    Span4Mux_h I__5889 (
            .O(N__25840),
            .I(N__25828));
    Span4Mux_s3_h I__5888 (
            .O(N__25837),
            .I(N__25823));
    LocalMux I__5887 (
            .O(N__25834),
            .I(N__25823));
    LocalMux I__5886 (
            .O(N__25831),
            .I(\Lab_UT.di_AMtens_2 ));
    Odrv4 I__5885 (
            .O(N__25828),
            .I(\Lab_UT.di_AMtens_2 ));
    Odrv4 I__5884 (
            .O(N__25823),
            .I(\Lab_UT.di_AMtens_2 ));
    InMux I__5883 (
            .O(N__25816),
            .I(N__25813));
    LocalMux I__5882 (
            .O(N__25813),
            .I(\Lab_UT.display.N_115 ));
    InMux I__5881 (
            .O(N__25810),
            .I(N__25806));
    CascadeMux I__5880 (
            .O(N__25809),
            .I(N__25803));
    LocalMux I__5879 (
            .O(N__25806),
            .I(N__25799));
    InMux I__5878 (
            .O(N__25803),
            .I(N__25796));
    InMux I__5877 (
            .O(N__25802),
            .I(N__25793));
    Span4Mux_s3_h I__5876 (
            .O(N__25799),
            .I(N__25788));
    LocalMux I__5875 (
            .O(N__25796),
            .I(N__25788));
    LocalMux I__5874 (
            .O(N__25793),
            .I(\Lab_UT.di_AStens_1 ));
    Odrv4 I__5873 (
            .O(N__25788),
            .I(\Lab_UT.di_AStens_1 ));
    CascadeMux I__5872 (
            .O(N__25783),
            .I(\Lab_UT.display.N_108_cascade_ ));
    InMux I__5871 (
            .O(N__25780),
            .I(N__25776));
    InMux I__5870 (
            .O(N__25779),
            .I(N__25772));
    LocalMux I__5869 (
            .O(N__25776),
            .I(N__25769));
    InMux I__5868 (
            .O(N__25775),
            .I(N__25766));
    LocalMux I__5867 (
            .O(N__25772),
            .I(N__25763));
    Span4Mux_v I__5866 (
            .O(N__25769),
            .I(N__25760));
    LocalMux I__5865 (
            .O(N__25766),
            .I(\Lab_UT.di_AMones_1 ));
    Odrv4 I__5864 (
            .O(N__25763),
            .I(\Lab_UT.di_AMones_1 ));
    Odrv4 I__5863 (
            .O(N__25760),
            .I(\Lab_UT.di_AMones_1 ));
    InMux I__5862 (
            .O(N__25753),
            .I(N__25750));
    LocalMux I__5861 (
            .O(N__25750),
            .I(N__25747));
    Span4Mux_h I__5860 (
            .O(N__25747),
            .I(N__25744));
    Odrv4 I__5859 (
            .O(N__25744),
            .I(\Lab_UT.display.dOutP_0_iv_i_0_1 ));
    CascadeMux I__5858 (
            .O(N__25741),
            .I(N__25738));
    InMux I__5857 (
            .O(N__25738),
            .I(N__25735));
    LocalMux I__5856 (
            .O(N__25735),
            .I(\Lab_UT.displayAlarmZ0Z_0 ));
    InMux I__5855 (
            .O(N__25732),
            .I(N__25729));
    LocalMux I__5854 (
            .O(N__25729),
            .I(N__25725));
    InMux I__5853 (
            .O(N__25728),
            .I(N__25721));
    Span4Mux_v I__5852 (
            .O(N__25725),
            .I(N__25718));
    InMux I__5851 (
            .O(N__25724),
            .I(N__25715));
    LocalMux I__5850 (
            .O(N__25721),
            .I(\Lab_UT.di_AStens_0 ));
    Odrv4 I__5849 (
            .O(N__25718),
            .I(\Lab_UT.di_AStens_0 ));
    LocalMux I__5848 (
            .O(N__25715),
            .I(\Lab_UT.di_AStens_0 ));
    InMux I__5847 (
            .O(N__25708),
            .I(N__25705));
    LocalMux I__5846 (
            .O(N__25705),
            .I(\Lab_UT.display.N_130 ));
    CascadeMux I__5845 (
            .O(N__25702),
            .I(\Lab_UT.display.dOutP_0_iv_i_0_0_cascade_ ));
    InMux I__5844 (
            .O(N__25699),
            .I(N__25696));
    LocalMux I__5843 (
            .O(N__25696),
            .I(N__25693));
    Span4Mux_v I__5842 (
            .O(N__25693),
            .I(N__25690));
    Odrv4 I__5841 (
            .O(N__25690),
            .I(\Lab_UT.display.dOutP_0_iv_i_1_0 ));
    CascadeMux I__5840 (
            .O(N__25687),
            .I(N__25684));
    InMux I__5839 (
            .O(N__25684),
            .I(N__25677));
    InMux I__5838 (
            .O(N__25683),
            .I(N__25677));
    InMux I__5837 (
            .O(N__25682),
            .I(N__25674));
    LocalMux I__5836 (
            .O(N__25677),
            .I(N__25671));
    LocalMux I__5835 (
            .O(N__25674),
            .I(N__25668));
    Span4Mux_h I__5834 (
            .O(N__25671),
            .I(N__25665));
    Odrv12 I__5833 (
            .O(N__25668),
            .I(L3_tx_data_0));
    Odrv4 I__5832 (
            .O(N__25665),
            .I(L3_tx_data_0));
    InMux I__5831 (
            .O(N__25660),
            .I(N__25654));
    InMux I__5830 (
            .O(N__25659),
            .I(N__25654));
    LocalMux I__5829 (
            .O(N__25654),
            .I(N__25651));
    Span4Mux_s2_h I__5828 (
            .O(N__25651),
            .I(N__25648));
    Odrv4 I__5827 (
            .O(N__25648),
            .I(\Lab_UT.display.N_153 ));
    CascadeMux I__5826 (
            .O(N__25645),
            .I(N__25642));
    InMux I__5825 (
            .O(N__25642),
            .I(N__25639));
    LocalMux I__5824 (
            .O(N__25639),
            .I(N__25636));
    Odrv4 I__5823 (
            .O(N__25636),
            .I(\Lab_UT.displayAlarmZ1Z_2 ));
    InMux I__5822 (
            .O(N__25633),
            .I(N__25630));
    LocalMux I__5821 (
            .O(N__25630),
            .I(N__25626));
    InMux I__5820 (
            .O(N__25629),
            .I(N__25622));
    Span4Mux_s2_h I__5819 (
            .O(N__25626),
            .I(N__25619));
    InMux I__5818 (
            .O(N__25625),
            .I(N__25616));
    LocalMux I__5817 (
            .O(N__25622),
            .I(\Lab_UT.di_AStens_2 ));
    Odrv4 I__5816 (
            .O(N__25619),
            .I(\Lab_UT.di_AStens_2 ));
    LocalMux I__5815 (
            .O(N__25616),
            .I(\Lab_UT.di_AStens_2 ));
    CascadeMux I__5814 (
            .O(N__25609),
            .I(\Lab_UT.display.dOutP_0_iv_i_0_2_cascade_ ));
    InMux I__5813 (
            .O(N__25606),
            .I(N__25603));
    LocalMux I__5812 (
            .O(N__25603),
            .I(N__25600));
    Span4Mux_v I__5811 (
            .O(N__25600),
            .I(N__25597));
    Odrv4 I__5810 (
            .O(N__25597),
            .I(\Lab_UT.display.dOutP_0_iv_i_1_2 ));
    CascadeMux I__5809 (
            .O(N__25594),
            .I(N__25591));
    InMux I__5808 (
            .O(N__25591),
            .I(N__25587));
    InMux I__5807 (
            .O(N__25590),
            .I(N__25583));
    LocalMux I__5806 (
            .O(N__25587),
            .I(N__25580));
    InMux I__5805 (
            .O(N__25586),
            .I(N__25577));
    LocalMux I__5804 (
            .O(N__25583),
            .I(N__25570));
    Span4Mux_s3_v I__5803 (
            .O(N__25580),
            .I(N__25570));
    LocalMux I__5802 (
            .O(N__25577),
            .I(N__25570));
    Odrv4 I__5801 (
            .O(N__25570),
            .I(L3_tx_data_2));
    InMux I__5800 (
            .O(N__25567),
            .I(N__25558));
    InMux I__5799 (
            .O(N__25566),
            .I(N__25558));
    InMux I__5798 (
            .O(N__25565),
            .I(N__25558));
    LocalMux I__5797 (
            .O(N__25558),
            .I(N__25555));
    Odrv4 I__5796 (
            .O(N__25555),
            .I(\Lab_UT.display.un42_dOutP_1 ));
    InMux I__5795 (
            .O(N__25552),
            .I(N__25546));
    InMux I__5794 (
            .O(N__25551),
            .I(N__25546));
    LocalMux I__5793 (
            .O(N__25546),
            .I(N__25543));
    Span4Mux_v I__5792 (
            .O(N__25543),
            .I(N__25540));
    Odrv4 I__5791 (
            .O(N__25540),
            .I(\Lab_UT.display.cnt_RNI1STE1Z0Z_1 ));
    CascadeMux I__5790 (
            .O(N__25537),
            .I(\Lab_UT.display.N_151_cascade_ ));
    InMux I__5789 (
            .O(N__25534),
            .I(N__25530));
    InMux I__5788 (
            .O(N__25533),
            .I(N__25527));
    LocalMux I__5787 (
            .O(N__25530),
            .I(N__25523));
    LocalMux I__5786 (
            .O(N__25527),
            .I(N__25520));
    InMux I__5785 (
            .O(N__25526),
            .I(N__25517));
    Span4Mux_s2_h I__5784 (
            .O(N__25523),
            .I(N__25514));
    Span4Mux_h I__5783 (
            .O(N__25520),
            .I(N__25511));
    LocalMux I__5782 (
            .O(N__25517),
            .I(\Lab_UT.di_AMtens_3 ));
    Odrv4 I__5781 (
            .O(N__25514),
            .I(\Lab_UT.di_AMtens_3 ));
    Odrv4 I__5780 (
            .O(N__25511),
            .I(\Lab_UT.di_AMtens_3 ));
    InMux I__5779 (
            .O(N__25504),
            .I(N__25501));
    LocalMux I__5778 (
            .O(N__25501),
            .I(N__25498));
    Odrv4 I__5777 (
            .O(N__25498),
            .I(\Lab_UT.display.N_124 ));
    CascadeMux I__5776 (
            .O(N__25495),
            .I(\Lab_UT.dictrl.decoder.de_littleNZ0Z_1_cascade_ ));
    InMux I__5775 (
            .O(N__25492),
            .I(N__25486));
    InMux I__5774 (
            .O(N__25491),
            .I(N__25479));
    InMux I__5773 (
            .O(N__25490),
            .I(N__25479));
    InMux I__5772 (
            .O(N__25489),
            .I(N__25479));
    LocalMux I__5771 (
            .O(N__25486),
            .I(N__25474));
    LocalMux I__5770 (
            .O(N__25479),
            .I(N__25471));
    InMux I__5769 (
            .O(N__25478),
            .I(N__25466));
    InMux I__5768 (
            .O(N__25477),
            .I(N__25466));
    Span4Mux_v I__5767 (
            .O(N__25474),
            .I(N__25461));
    Span4Mux_v I__5766 (
            .O(N__25471),
            .I(N__25461));
    LocalMux I__5765 (
            .O(N__25466),
            .I(Lab_UT_dictrl_decoder_de_cr_2));
    Odrv4 I__5764 (
            .O(N__25461),
            .I(Lab_UT_dictrl_decoder_de_cr_2));
    CascadeMux I__5763 (
            .O(N__25456),
            .I(N__25453));
    InMux I__5762 (
            .O(N__25453),
            .I(N__25447));
    InMux I__5761 (
            .O(N__25452),
            .I(N__25447));
    LocalMux I__5760 (
            .O(N__25447),
            .I(N__25444));
    Span4Mux_v I__5759 (
            .O(N__25444),
            .I(N__25441));
    Span4Mux_v I__5758 (
            .O(N__25441),
            .I(N__25438));
    Odrv4 I__5757 (
            .O(N__25438),
            .I(\Lab_UT.n_rdy ));
    InMux I__5756 (
            .O(N__25435),
            .I(N__25432));
    LocalMux I__5755 (
            .O(N__25432),
            .I(\resetGen.escKeyZ0Z_3 ));
    CEMux I__5754 (
            .O(N__25429),
            .I(N__25408));
    CEMux I__5753 (
            .O(N__25428),
            .I(N__25408));
    CEMux I__5752 (
            .O(N__25427),
            .I(N__25408));
    CEMux I__5751 (
            .O(N__25426),
            .I(N__25408));
    CEMux I__5750 (
            .O(N__25425),
            .I(N__25408));
    CEMux I__5749 (
            .O(N__25424),
            .I(N__25408));
    CEMux I__5748 (
            .O(N__25423),
            .I(N__25408));
    GlobalMux I__5747 (
            .O(N__25408),
            .I(N__25405));
    gio2CtrlBuf I__5746 (
            .O(N__25405),
            .I(\buart.Z_rx.sample_g ));
    InMux I__5745 (
            .O(N__25402),
            .I(N__25399));
    LocalMux I__5744 (
            .O(N__25399),
            .I(N__25391));
    InMux I__5743 (
            .O(N__25398),
            .I(N__25386));
    InMux I__5742 (
            .O(N__25397),
            .I(N__25386));
    InMux I__5741 (
            .O(N__25396),
            .I(N__25381));
    InMux I__5740 (
            .O(N__25395),
            .I(N__25381));
    InMux I__5739 (
            .O(N__25394),
            .I(N__25378));
    Span4Mux_s3_h I__5738 (
            .O(N__25391),
            .I(N__25363));
    LocalMux I__5737 (
            .O(N__25386),
            .I(N__25363));
    LocalMux I__5736 (
            .O(N__25381),
            .I(N__25363));
    LocalMux I__5735 (
            .O(N__25378),
            .I(N__25363));
    InMux I__5734 (
            .O(N__25377),
            .I(N__25360));
    InMux I__5733 (
            .O(N__25376),
            .I(N__25357));
    InMux I__5732 (
            .O(N__25375),
            .I(N__25350));
    InMux I__5731 (
            .O(N__25374),
            .I(N__25350));
    InMux I__5730 (
            .O(N__25373),
            .I(N__25350));
    InMux I__5729 (
            .O(N__25372),
            .I(N__25347));
    Span4Mux_h I__5728 (
            .O(N__25363),
            .I(N__25341));
    LocalMux I__5727 (
            .O(N__25360),
            .I(N__25334));
    LocalMux I__5726 (
            .O(N__25357),
            .I(N__25334));
    LocalMux I__5725 (
            .O(N__25350),
            .I(N__25334));
    LocalMux I__5724 (
            .O(N__25347),
            .I(N__25331));
    InMux I__5723 (
            .O(N__25346),
            .I(N__25324));
    InMux I__5722 (
            .O(N__25345),
            .I(N__25324));
    InMux I__5721 (
            .O(N__25344),
            .I(N__25324));
    Odrv4 I__5720 (
            .O(N__25341),
            .I(bu_rx_data_7));
    Odrv12 I__5719 (
            .O(N__25334),
            .I(bu_rx_data_7));
    Odrv4 I__5718 (
            .O(N__25331),
            .I(bu_rx_data_7));
    LocalMux I__5717 (
            .O(N__25324),
            .I(bu_rx_data_7));
    InMux I__5716 (
            .O(N__25315),
            .I(N__25308));
    InMux I__5715 (
            .O(N__25314),
            .I(N__25308));
    InMux I__5714 (
            .O(N__25313),
            .I(N__25305));
    LocalMux I__5713 (
            .O(N__25308),
            .I(N__25297));
    LocalMux I__5712 (
            .O(N__25305),
            .I(N__25294));
    InMux I__5711 (
            .O(N__25304),
            .I(N__25291));
    InMux I__5710 (
            .O(N__25303),
            .I(N__25288));
    InMux I__5709 (
            .O(N__25302),
            .I(N__25283));
    InMux I__5708 (
            .O(N__25301),
            .I(N__25283));
    InMux I__5707 (
            .O(N__25300),
            .I(N__25280));
    Span4Mux_v I__5706 (
            .O(N__25297),
            .I(N__25274));
    Span4Mux_s2_v I__5705 (
            .O(N__25294),
            .I(N__25274));
    LocalMux I__5704 (
            .O(N__25291),
            .I(N__25269));
    LocalMux I__5703 (
            .O(N__25288),
            .I(N__25266));
    LocalMux I__5702 (
            .O(N__25283),
            .I(N__25261));
    LocalMux I__5701 (
            .O(N__25280),
            .I(N__25261));
    InMux I__5700 (
            .O(N__25279),
            .I(N__25257));
    Span4Mux_h I__5699 (
            .O(N__25274),
            .I(N__25254));
    InMux I__5698 (
            .O(N__25273),
            .I(N__25251));
    InMux I__5697 (
            .O(N__25272),
            .I(N__25248));
    Span4Mux_v I__5696 (
            .O(N__25269),
            .I(N__25241));
    Span4Mux_h I__5695 (
            .O(N__25266),
            .I(N__25241));
    Span4Mux_s2_v I__5694 (
            .O(N__25261),
            .I(N__25241));
    InMux I__5693 (
            .O(N__25260),
            .I(N__25238));
    LocalMux I__5692 (
            .O(N__25257),
            .I(bu_rx_data_4));
    Odrv4 I__5691 (
            .O(N__25254),
            .I(bu_rx_data_4));
    LocalMux I__5690 (
            .O(N__25251),
            .I(bu_rx_data_4));
    LocalMux I__5689 (
            .O(N__25248),
            .I(bu_rx_data_4));
    Odrv4 I__5688 (
            .O(N__25241),
            .I(bu_rx_data_4));
    LocalMux I__5687 (
            .O(N__25238),
            .I(bu_rx_data_4));
    InMux I__5686 (
            .O(N__25225),
            .I(N__25222));
    LocalMux I__5685 (
            .O(N__25222),
            .I(N__25219));
    Odrv4 I__5684 (
            .O(N__25219),
            .I(\Lab_UT.dictrl.decoder.de_atSignZ0Z_5 ));
    CascadeMux I__5683 (
            .O(N__25216),
            .I(N__25213));
    InMux I__5682 (
            .O(N__25213),
            .I(N__25201));
    InMux I__5681 (
            .O(N__25212),
            .I(N__25201));
    InMux I__5680 (
            .O(N__25211),
            .I(N__25201));
    InMux I__5679 (
            .O(N__25210),
            .I(N__25201));
    LocalMux I__5678 (
            .O(N__25201),
            .I(N__25196));
    InMux I__5677 (
            .O(N__25200),
            .I(N__25193));
    InMux I__5676 (
            .O(N__25199),
            .I(N__25190));
    Sp12to4 I__5675 (
            .O(N__25196),
            .I(N__25185));
    LocalMux I__5674 (
            .O(N__25193),
            .I(N__25185));
    LocalMux I__5673 (
            .O(N__25190),
            .I(\Lab_UT.uu0.l_precountZ0Z_0 ));
    Odrv12 I__5672 (
            .O(N__25185),
            .I(\Lab_UT.uu0.l_precountZ0Z_0 ));
    InMux I__5671 (
            .O(N__25180),
            .I(N__25176));
    InMux I__5670 (
            .O(N__25179),
            .I(N__25173));
    LocalMux I__5669 (
            .O(N__25176),
            .I(N__25170));
    LocalMux I__5668 (
            .O(N__25173),
            .I(N__25167));
    Span4Mux_v I__5667 (
            .O(N__25170),
            .I(N__25162));
    Span4Mux_s2_h I__5666 (
            .O(N__25167),
            .I(N__25162));
    Span4Mux_h I__5665 (
            .O(N__25162),
            .I(N__25157));
    InMux I__5664 (
            .O(N__25161),
            .I(N__25152));
    InMux I__5663 (
            .O(N__25160),
            .I(N__25152));
    Odrv4 I__5662 (
            .O(N__25157),
            .I(\uu2.un404_ci_0 ));
    LocalMux I__5661 (
            .O(N__25152),
            .I(\uu2.un404_ci_0 ));
    InMux I__5660 (
            .O(N__25147),
            .I(N__25143));
    InMux I__5659 (
            .O(N__25146),
            .I(N__25140));
    LocalMux I__5658 (
            .O(N__25143),
            .I(N__25137));
    LocalMux I__5657 (
            .O(N__25140),
            .I(N__25134));
    Span4Mux_v I__5656 (
            .O(N__25137),
            .I(N__25126));
    Span4Mux_s3_h I__5655 (
            .O(N__25134),
            .I(N__25126));
    InMux I__5654 (
            .O(N__25133),
            .I(N__25119));
    InMux I__5653 (
            .O(N__25132),
            .I(N__25119));
    InMux I__5652 (
            .O(N__25131),
            .I(N__25119));
    Odrv4 I__5651 (
            .O(N__25126),
            .I(\uu2.trig_rd_is_det ));
    LocalMux I__5650 (
            .O(N__25119),
            .I(\uu2.trig_rd_is_det ));
    CascadeMux I__5649 (
            .O(N__25114),
            .I(N__25111));
    InMux I__5648 (
            .O(N__25111),
            .I(N__25105));
    InMux I__5647 (
            .O(N__25110),
            .I(N__25100));
    InMux I__5646 (
            .O(N__25109),
            .I(N__25100));
    InMux I__5645 (
            .O(N__25108),
            .I(N__25097));
    LocalMux I__5644 (
            .O(N__25105),
            .I(N__25092));
    LocalMux I__5643 (
            .O(N__25100),
            .I(N__25092));
    LocalMux I__5642 (
            .O(N__25097),
            .I(N__25089));
    Span4Mux_h I__5641 (
            .O(N__25092),
            .I(N__25085));
    Span4Mux_h I__5640 (
            .O(N__25089),
            .I(N__25082));
    InMux I__5639 (
            .O(N__25088),
            .I(N__25079));
    Span4Mux_h I__5638 (
            .O(N__25085),
            .I(N__25076));
    Odrv4 I__5637 (
            .O(N__25082),
            .I(\uu2.r_addrZ0Z_4 ));
    LocalMux I__5636 (
            .O(N__25079),
            .I(\uu2.r_addrZ0Z_4 ));
    Odrv4 I__5635 (
            .O(N__25076),
            .I(\uu2.r_addrZ0Z_4 ));
    InMux I__5634 (
            .O(N__25069),
            .I(N__25066));
    LocalMux I__5633 (
            .O(N__25066),
            .I(N__25063));
    Span12Mux_s8_v I__5632 (
            .O(N__25063),
            .I(N__25058));
    InMux I__5631 (
            .O(N__25062),
            .I(N__25053));
    InMux I__5630 (
            .O(N__25061),
            .I(N__25053));
    Odrv12 I__5629 (
            .O(N__25058),
            .I(\Lab_UT.di_AMtens_0 ));
    LocalMux I__5628 (
            .O(N__25053),
            .I(\Lab_UT.di_AMtens_0 ));
    CascadeMux I__5627 (
            .O(N__25048),
            .I(N__25042));
    CascadeMux I__5626 (
            .O(N__25047),
            .I(N__25036));
    CascadeMux I__5625 (
            .O(N__25046),
            .I(N__25033));
    InMux I__5624 (
            .O(N__25045),
            .I(N__25026));
    InMux I__5623 (
            .O(N__25042),
            .I(N__25026));
    InMux I__5622 (
            .O(N__25041),
            .I(N__25026));
    InMux I__5621 (
            .O(N__25040),
            .I(N__25016));
    CascadeMux I__5620 (
            .O(N__25039),
            .I(N__25013));
    InMux I__5619 (
            .O(N__25036),
            .I(N__25005));
    InMux I__5618 (
            .O(N__25033),
            .I(N__25002));
    LocalMux I__5617 (
            .O(N__25026),
            .I(N__24999));
    InMux I__5616 (
            .O(N__25025),
            .I(N__24996));
    InMux I__5615 (
            .O(N__25024),
            .I(N__24987));
    InMux I__5614 (
            .O(N__25023),
            .I(N__24987));
    InMux I__5613 (
            .O(N__25022),
            .I(N__24987));
    InMux I__5612 (
            .O(N__25021),
            .I(N__24987));
    InMux I__5611 (
            .O(N__25020),
            .I(N__24982));
    InMux I__5610 (
            .O(N__25019),
            .I(N__24982));
    LocalMux I__5609 (
            .O(N__25016),
            .I(N__24979));
    InMux I__5608 (
            .O(N__25013),
            .I(N__24976));
    InMux I__5607 (
            .O(N__25012),
            .I(N__24973));
    InMux I__5606 (
            .O(N__25011),
            .I(N__24968));
    InMux I__5605 (
            .O(N__25010),
            .I(N__24968));
    CascadeMux I__5604 (
            .O(N__25009),
            .I(N__24965));
    InMux I__5603 (
            .O(N__25008),
            .I(N__24961));
    LocalMux I__5602 (
            .O(N__25005),
            .I(N__24958));
    LocalMux I__5601 (
            .O(N__25002),
            .I(N__24953));
    Span4Mux_s2_h I__5600 (
            .O(N__24999),
            .I(N__24953));
    LocalMux I__5599 (
            .O(N__24996),
            .I(N__24950));
    LocalMux I__5598 (
            .O(N__24987),
            .I(N__24947));
    LocalMux I__5597 (
            .O(N__24982),
            .I(N__24944));
    Span4Mux_h I__5596 (
            .O(N__24979),
            .I(N__24935));
    LocalMux I__5595 (
            .O(N__24976),
            .I(N__24935));
    LocalMux I__5594 (
            .O(N__24973),
            .I(N__24935));
    LocalMux I__5593 (
            .O(N__24968),
            .I(N__24935));
    InMux I__5592 (
            .O(N__24965),
            .I(N__24930));
    InMux I__5591 (
            .O(N__24964),
            .I(N__24930));
    LocalMux I__5590 (
            .O(N__24961),
            .I(N__24927));
    Span4Mux_h I__5589 (
            .O(N__24958),
            .I(N__24922));
    Span4Mux_h I__5588 (
            .O(N__24953),
            .I(N__24922));
    Span4Mux_v I__5587 (
            .O(N__24950),
            .I(N__24919));
    Span4Mux_v I__5586 (
            .O(N__24947),
            .I(N__24910));
    Span4Mux_h I__5585 (
            .O(N__24944),
            .I(N__24910));
    Span4Mux_v I__5584 (
            .O(N__24935),
            .I(N__24910));
    LocalMux I__5583 (
            .O(N__24930),
            .I(N__24910));
    Odrv12 I__5582 (
            .O(N__24927),
            .I(\Lab_UT.dictrl.currStateZ0Z_2 ));
    Odrv4 I__5581 (
            .O(N__24922),
            .I(\Lab_UT.dictrl.currStateZ0Z_2 ));
    Odrv4 I__5580 (
            .O(N__24919),
            .I(\Lab_UT.dictrl.currStateZ0Z_2 ));
    Odrv4 I__5579 (
            .O(N__24910),
            .I(\Lab_UT.dictrl.currStateZ0Z_2 ));
    CascadeMux I__5578 (
            .O(N__24901),
            .I(N__24894));
    CascadeMux I__5577 (
            .O(N__24900),
            .I(N__24891));
    CascadeMux I__5576 (
            .O(N__24899),
            .I(N__24882));
    CascadeMux I__5575 (
            .O(N__24898),
            .I(N__24879));
    CascadeMux I__5574 (
            .O(N__24897),
            .I(N__24875));
    InMux I__5573 (
            .O(N__24894),
            .I(N__24871));
    InMux I__5572 (
            .O(N__24891),
            .I(N__24868));
    InMux I__5571 (
            .O(N__24890),
            .I(N__24865));
    InMux I__5570 (
            .O(N__24889),
            .I(N__24856));
    InMux I__5569 (
            .O(N__24888),
            .I(N__24856));
    InMux I__5568 (
            .O(N__24887),
            .I(N__24849));
    InMux I__5567 (
            .O(N__24886),
            .I(N__24849));
    InMux I__5566 (
            .O(N__24885),
            .I(N__24849));
    InMux I__5565 (
            .O(N__24882),
            .I(N__24844));
    InMux I__5564 (
            .O(N__24879),
            .I(N__24844));
    InMux I__5563 (
            .O(N__24878),
            .I(N__24841));
    InMux I__5562 (
            .O(N__24875),
            .I(N__24838));
    InMux I__5561 (
            .O(N__24874),
            .I(N__24835));
    LocalMux I__5560 (
            .O(N__24871),
            .I(N__24830));
    LocalMux I__5559 (
            .O(N__24868),
            .I(N__24830));
    LocalMux I__5558 (
            .O(N__24865),
            .I(N__24827));
    InMux I__5557 (
            .O(N__24864),
            .I(N__24824));
    InMux I__5556 (
            .O(N__24863),
            .I(N__24819));
    InMux I__5555 (
            .O(N__24862),
            .I(N__24819));
    CascadeMux I__5554 (
            .O(N__24861),
            .I(N__24816));
    LocalMux I__5553 (
            .O(N__24856),
            .I(N__24810));
    LocalMux I__5552 (
            .O(N__24849),
            .I(N__24807));
    LocalMux I__5551 (
            .O(N__24844),
            .I(N__24804));
    LocalMux I__5550 (
            .O(N__24841),
            .I(N__24797));
    LocalMux I__5549 (
            .O(N__24838),
            .I(N__24797));
    LocalMux I__5548 (
            .O(N__24835),
            .I(N__24790));
    Span4Mux_s3_h I__5547 (
            .O(N__24830),
            .I(N__24790));
    Span4Mux_h I__5546 (
            .O(N__24827),
            .I(N__24790));
    LocalMux I__5545 (
            .O(N__24824),
            .I(N__24787));
    LocalMux I__5544 (
            .O(N__24819),
            .I(N__24784));
    InMux I__5543 (
            .O(N__24816),
            .I(N__24779));
    InMux I__5542 (
            .O(N__24815),
            .I(N__24779));
    InMux I__5541 (
            .O(N__24814),
            .I(N__24774));
    InMux I__5540 (
            .O(N__24813),
            .I(N__24774));
    Span4Mux_v I__5539 (
            .O(N__24810),
            .I(N__24767));
    Span4Mux_h I__5538 (
            .O(N__24807),
            .I(N__24767));
    Span4Mux_v I__5537 (
            .O(N__24804),
            .I(N__24767));
    InMux I__5536 (
            .O(N__24803),
            .I(N__24762));
    InMux I__5535 (
            .O(N__24802),
            .I(N__24762));
    Span4Mux_s3_h I__5534 (
            .O(N__24797),
            .I(N__24757));
    Span4Mux_h I__5533 (
            .O(N__24790),
            .I(N__24757));
    Odrv4 I__5532 (
            .O(N__24787),
            .I(\Lab_UT.dictrl.currState_i_5_3 ));
    Odrv4 I__5531 (
            .O(N__24784),
            .I(\Lab_UT.dictrl.currState_i_5_3 ));
    LocalMux I__5530 (
            .O(N__24779),
            .I(\Lab_UT.dictrl.currState_i_5_3 ));
    LocalMux I__5529 (
            .O(N__24774),
            .I(\Lab_UT.dictrl.currState_i_5_3 ));
    Odrv4 I__5528 (
            .O(N__24767),
            .I(\Lab_UT.dictrl.currState_i_5_3 ));
    LocalMux I__5527 (
            .O(N__24762),
            .I(\Lab_UT.dictrl.currState_i_5_3 ));
    Odrv4 I__5526 (
            .O(N__24757),
            .I(\Lab_UT.dictrl.currState_i_5_3 ));
    CascadeMux I__5525 (
            .O(N__24742),
            .I(N__24739));
    InMux I__5524 (
            .O(N__24739),
            .I(N__24736));
    LocalMux I__5523 (
            .O(N__24736),
            .I(N__24733));
    Odrv4 I__5522 (
            .O(N__24733),
            .I(\Lab_UT.dictrl.r_dicRun_r_1 ));
    CascadeMux I__5521 (
            .O(N__24730),
            .I(N__24727));
    InMux I__5520 (
            .O(N__24727),
            .I(N__24720));
    InMux I__5519 (
            .O(N__24726),
            .I(N__24720));
    InMux I__5518 (
            .O(N__24725),
            .I(N__24717));
    LocalMux I__5517 (
            .O(N__24720),
            .I(N__24714));
    LocalMux I__5516 (
            .O(N__24717),
            .I(N__24711));
    Odrv4 I__5515 (
            .O(N__24714),
            .I(\Lab_UT.dictrl.r_dicLdMtens15_1i ));
    Odrv4 I__5514 (
            .O(N__24711),
            .I(\Lab_UT.dictrl.r_dicLdMtens15_1i ));
    InMux I__5513 (
            .O(N__24706),
            .I(N__24699));
    InMux I__5512 (
            .O(N__24705),
            .I(N__24696));
    InMux I__5511 (
            .O(N__24704),
            .I(N__24690));
    InMux I__5510 (
            .O(N__24703),
            .I(N__24690));
    IoInMux I__5509 (
            .O(N__24702),
            .I(N__24666));
    LocalMux I__5508 (
            .O(N__24699),
            .I(N__24663));
    LocalMux I__5507 (
            .O(N__24696),
            .I(N__24660));
    InMux I__5506 (
            .O(N__24695),
            .I(N__24657));
    LocalMux I__5505 (
            .O(N__24690),
            .I(N__24654));
    InMux I__5504 (
            .O(N__24689),
            .I(N__24651));
    InMux I__5503 (
            .O(N__24688),
            .I(N__24644));
    InMux I__5502 (
            .O(N__24687),
            .I(N__24644));
    InMux I__5501 (
            .O(N__24686),
            .I(N__24644));
    InMux I__5500 (
            .O(N__24685),
            .I(N__24637));
    InMux I__5499 (
            .O(N__24684),
            .I(N__24637));
    InMux I__5498 (
            .O(N__24683),
            .I(N__24637));
    InMux I__5497 (
            .O(N__24682),
            .I(N__24634));
    InMux I__5496 (
            .O(N__24681),
            .I(N__24631));
    InMux I__5495 (
            .O(N__24680),
            .I(N__24628));
    InMux I__5494 (
            .O(N__24679),
            .I(N__24623));
    InMux I__5493 (
            .O(N__24678),
            .I(N__24618));
    InMux I__5492 (
            .O(N__24677),
            .I(N__24618));
    InMux I__5491 (
            .O(N__24676),
            .I(N__24615));
    InMux I__5490 (
            .O(N__24675),
            .I(N__24606));
    InMux I__5489 (
            .O(N__24674),
            .I(N__24606));
    InMux I__5488 (
            .O(N__24673),
            .I(N__24606));
    InMux I__5487 (
            .O(N__24672),
            .I(N__24606));
    InMux I__5486 (
            .O(N__24671),
            .I(N__24599));
    InMux I__5485 (
            .O(N__24670),
            .I(N__24599));
    InMux I__5484 (
            .O(N__24669),
            .I(N__24599));
    LocalMux I__5483 (
            .O(N__24666),
            .I(N__24596));
    Span4Mux_v I__5482 (
            .O(N__24663),
            .I(N__24591));
    Span4Mux_v I__5481 (
            .O(N__24660),
            .I(N__24591));
    LocalMux I__5480 (
            .O(N__24657),
            .I(N__24584));
    Span4Mux_s3_v I__5479 (
            .O(N__24654),
            .I(N__24584));
    LocalMux I__5478 (
            .O(N__24651),
            .I(N__24584));
    LocalMux I__5477 (
            .O(N__24644),
            .I(N__24579));
    LocalMux I__5476 (
            .O(N__24637),
            .I(N__24579));
    LocalMux I__5475 (
            .O(N__24634),
            .I(N__24574));
    LocalMux I__5474 (
            .O(N__24631),
            .I(N__24569));
    LocalMux I__5473 (
            .O(N__24628),
            .I(N__24569));
    InMux I__5472 (
            .O(N__24627),
            .I(N__24564));
    InMux I__5471 (
            .O(N__24626),
            .I(N__24564));
    LocalMux I__5470 (
            .O(N__24623),
            .I(N__24557));
    LocalMux I__5469 (
            .O(N__24618),
            .I(N__24557));
    LocalMux I__5468 (
            .O(N__24615),
            .I(N__24557));
    LocalMux I__5467 (
            .O(N__24606),
            .I(N__24550));
    LocalMux I__5466 (
            .O(N__24599),
            .I(N__24550));
    IoSpan4Mux I__5465 (
            .O(N__24596),
            .I(N__24550));
    Span4Mux_h I__5464 (
            .O(N__24591),
            .I(N__24547));
    Span4Mux_v I__5463 (
            .O(N__24584),
            .I(N__24542));
    Span4Mux_v I__5462 (
            .O(N__24579),
            .I(N__24542));
    InMux I__5461 (
            .O(N__24578),
            .I(N__24537));
    InMux I__5460 (
            .O(N__24577),
            .I(N__24537));
    Span4Mux_h I__5459 (
            .O(N__24574),
            .I(N__24532));
    Span4Mux_s3_h I__5458 (
            .O(N__24569),
            .I(N__24532));
    LocalMux I__5457 (
            .O(N__24564),
            .I(N__24525));
    Span4Mux_h I__5456 (
            .O(N__24557),
            .I(N__24525));
    Span4Mux_s3_h I__5455 (
            .O(N__24550),
            .I(N__24525));
    Odrv4 I__5454 (
            .O(N__24547),
            .I(rst));
    Odrv4 I__5453 (
            .O(N__24542),
            .I(rst));
    LocalMux I__5452 (
            .O(N__24537),
            .I(rst));
    Odrv4 I__5451 (
            .O(N__24532),
            .I(rst));
    Odrv4 I__5450 (
            .O(N__24525),
            .I(rst));
    InMux I__5449 (
            .O(N__24514),
            .I(N__24509));
    InMux I__5448 (
            .O(N__24513),
            .I(N__24504));
    InMux I__5447 (
            .O(N__24512),
            .I(N__24504));
    LocalMux I__5446 (
            .O(N__24509),
            .I(\Lab_UT.dictrl.r_dicLdMtens15_1 ));
    LocalMux I__5445 (
            .O(N__24504),
            .I(\Lab_UT.dictrl.r_dicLdMtens15_1 ));
    CascadeMux I__5444 (
            .O(N__24499),
            .I(\Lab_UT.dictrl.decoder.de_atSignZ0Z_4_cascade_ ));
    InMux I__5443 (
            .O(N__24496),
            .I(N__24490));
    InMux I__5442 (
            .O(N__24495),
            .I(N__24490));
    LocalMux I__5441 (
            .O(N__24490),
            .I(N__24487));
    Odrv4 I__5440 (
            .O(N__24487),
            .I(\Lab_UT.dictrl.de_atSign ));
    CascadeMux I__5439 (
            .O(N__24484),
            .I(\Lab_UT.dictrl.de_littleA_2_cascade_ ));
    InMux I__5438 (
            .O(N__24481),
            .I(N__24478));
    LocalMux I__5437 (
            .O(N__24478),
            .I(N__24472));
    InMux I__5436 (
            .O(N__24477),
            .I(N__24469));
    InMux I__5435 (
            .O(N__24476),
            .I(N__24466));
    InMux I__5434 (
            .O(N__24475),
            .I(N__24463));
    Span4Mux_h I__5433 (
            .O(N__24472),
            .I(N__24460));
    LocalMux I__5432 (
            .O(N__24469),
            .I(N__24457));
    LocalMux I__5431 (
            .O(N__24466),
            .I(\Lab_UT.dictrl.de_littleL ));
    LocalMux I__5430 (
            .O(N__24463),
            .I(\Lab_UT.dictrl.de_littleL ));
    Odrv4 I__5429 (
            .O(N__24460),
            .I(\Lab_UT.dictrl.de_littleL ));
    Odrv12 I__5428 (
            .O(N__24457),
            .I(\Lab_UT.dictrl.de_littleL ));
    InMux I__5427 (
            .O(N__24448),
            .I(N__24437));
    InMux I__5426 (
            .O(N__24447),
            .I(N__24434));
    InMux I__5425 (
            .O(N__24446),
            .I(N__24429));
    InMux I__5424 (
            .O(N__24445),
            .I(N__24429));
    InMux I__5423 (
            .O(N__24444),
            .I(N__24426));
    InMux I__5422 (
            .O(N__24443),
            .I(N__24423));
    InMux I__5421 (
            .O(N__24442),
            .I(N__24418));
    InMux I__5420 (
            .O(N__24441),
            .I(N__24418));
    InMux I__5419 (
            .O(N__24440),
            .I(N__24411));
    LocalMux I__5418 (
            .O(N__24437),
            .I(N__24408));
    LocalMux I__5417 (
            .O(N__24434),
            .I(N__24401));
    LocalMux I__5416 (
            .O(N__24429),
            .I(N__24401));
    LocalMux I__5415 (
            .O(N__24426),
            .I(N__24401));
    LocalMux I__5414 (
            .O(N__24423),
            .I(N__24398));
    LocalMux I__5413 (
            .O(N__24418),
            .I(N__24395));
    InMux I__5412 (
            .O(N__24417),
            .I(N__24392));
    InMux I__5411 (
            .O(N__24416),
            .I(N__24387));
    InMux I__5410 (
            .O(N__24415),
            .I(N__24387));
    InMux I__5409 (
            .O(N__24414),
            .I(N__24384));
    LocalMux I__5408 (
            .O(N__24411),
            .I(N__24379));
    Span4Mux_v I__5407 (
            .O(N__24408),
            .I(N__24379));
    Span4Mux_h I__5406 (
            .O(N__24401),
            .I(N__24376));
    Span4Mux_h I__5405 (
            .O(N__24398),
            .I(N__24371));
    Span4Mux_s2_v I__5404 (
            .O(N__24395),
            .I(N__24371));
    LocalMux I__5403 (
            .O(N__24392),
            .I(bu_rx_data_5));
    LocalMux I__5402 (
            .O(N__24387),
            .I(bu_rx_data_5));
    LocalMux I__5401 (
            .O(N__24384),
            .I(bu_rx_data_5));
    Odrv4 I__5400 (
            .O(N__24379),
            .I(bu_rx_data_5));
    Odrv4 I__5399 (
            .O(N__24376),
            .I(bu_rx_data_5));
    Odrv4 I__5398 (
            .O(N__24371),
            .I(bu_rx_data_5));
    InMux I__5397 (
            .O(N__24358),
            .I(N__24351));
    InMux I__5396 (
            .O(N__24357),
            .I(N__24351));
    InMux I__5395 (
            .O(N__24356),
            .I(N__24348));
    LocalMux I__5394 (
            .O(N__24351),
            .I(N__24344));
    LocalMux I__5393 (
            .O(N__24348),
            .I(N__24341));
    InMux I__5392 (
            .O(N__24347),
            .I(N__24337));
    Span4Mux_v I__5391 (
            .O(N__24344),
            .I(N__24332));
    Span4Mux_s2_v I__5390 (
            .O(N__24341),
            .I(N__24332));
    InMux I__5389 (
            .O(N__24340),
            .I(N__24329));
    LocalMux I__5388 (
            .O(N__24337),
            .I(\Lab_UT.dictrl.de_littleL_4 ));
    Odrv4 I__5387 (
            .O(N__24332),
            .I(\Lab_UT.dictrl.de_littleL_4 ));
    LocalMux I__5386 (
            .O(N__24329),
            .I(\Lab_UT.dictrl.de_littleL_4 ));
    CascadeMux I__5385 (
            .O(N__24322),
            .I(N__24317));
    CascadeMux I__5384 (
            .O(N__24321),
            .I(N__24314));
    CascadeMux I__5383 (
            .O(N__24320),
            .I(N__24311));
    InMux I__5382 (
            .O(N__24317),
            .I(N__24301));
    InMux I__5381 (
            .O(N__24314),
            .I(N__24301));
    InMux I__5380 (
            .O(N__24311),
            .I(N__24301));
    CascadeMux I__5379 (
            .O(N__24310),
            .I(N__24297));
    InMux I__5378 (
            .O(N__24309),
            .I(N__24291));
    InMux I__5377 (
            .O(N__24308),
            .I(N__24288));
    LocalMux I__5376 (
            .O(N__24301),
            .I(N__24285));
    InMux I__5375 (
            .O(N__24300),
            .I(N__24282));
    InMux I__5374 (
            .O(N__24297),
            .I(N__24275));
    InMux I__5373 (
            .O(N__24296),
            .I(N__24275));
    InMux I__5372 (
            .O(N__24295),
            .I(N__24275));
    CascadeMux I__5371 (
            .O(N__24294),
            .I(N__24272));
    LocalMux I__5370 (
            .O(N__24291),
            .I(N__24267));
    LocalMux I__5369 (
            .O(N__24288),
            .I(N__24263));
    Span4Mux_s3_h I__5368 (
            .O(N__24285),
            .I(N__24260));
    LocalMux I__5367 (
            .O(N__24282),
            .I(N__24255));
    LocalMux I__5366 (
            .O(N__24275),
            .I(N__24255));
    InMux I__5365 (
            .O(N__24272),
            .I(N__24252));
    InMux I__5364 (
            .O(N__24271),
            .I(N__24247));
    InMux I__5363 (
            .O(N__24270),
            .I(N__24247));
    Span4Mux_v I__5362 (
            .O(N__24267),
            .I(N__24244));
    InMux I__5361 (
            .O(N__24266),
            .I(N__24241));
    Span4Mux_h I__5360 (
            .O(N__24263),
            .I(N__24238));
    Span4Mux_h I__5359 (
            .O(N__24260),
            .I(N__24235));
    Span4Mux_v I__5358 (
            .O(N__24255),
            .I(N__24230));
    LocalMux I__5357 (
            .O(N__24252),
            .I(N__24230));
    LocalMux I__5356 (
            .O(N__24247),
            .I(bu_rx_data_6));
    Odrv4 I__5355 (
            .O(N__24244),
            .I(bu_rx_data_6));
    LocalMux I__5354 (
            .O(N__24241),
            .I(bu_rx_data_6));
    Odrv4 I__5353 (
            .O(N__24238),
            .I(bu_rx_data_6));
    Odrv4 I__5352 (
            .O(N__24235),
            .I(bu_rx_data_6));
    Odrv4 I__5351 (
            .O(N__24230),
            .I(bu_rx_data_6));
    InMux I__5350 (
            .O(N__24217),
            .I(N__24214));
    LocalMux I__5349 (
            .O(N__24214),
            .I(N__24211));
    Odrv4 I__5348 (
            .O(N__24211),
            .I(\Lab_UT.dictrl.g0_4_2 ));
    CascadeMux I__5347 (
            .O(N__24208),
            .I(N__24203));
    InMux I__5346 (
            .O(N__24207),
            .I(N__24200));
    CascadeMux I__5345 (
            .O(N__24206),
            .I(N__24197));
    InMux I__5344 (
            .O(N__24203),
            .I(N__24194));
    LocalMux I__5343 (
            .O(N__24200),
            .I(N__24191));
    InMux I__5342 (
            .O(N__24197),
            .I(N__24188));
    LocalMux I__5341 (
            .O(N__24194),
            .I(N__24185));
    Odrv12 I__5340 (
            .O(N__24191),
            .I(\Lab_UT.dictrl.de_littleA_2 ));
    LocalMux I__5339 (
            .O(N__24188),
            .I(\Lab_UT.dictrl.de_littleA_2 ));
    Odrv4 I__5338 (
            .O(N__24185),
            .I(\Lab_UT.dictrl.de_littleA_2 ));
    InMux I__5337 (
            .O(N__24178),
            .I(N__24173));
    CascadeMux I__5336 (
            .O(N__24177),
            .I(N__24169));
    CascadeMux I__5335 (
            .O(N__24176),
            .I(N__24165));
    LocalMux I__5334 (
            .O(N__24173),
            .I(N__24162));
    InMux I__5333 (
            .O(N__24172),
            .I(N__24159));
    InMux I__5332 (
            .O(N__24169),
            .I(N__24150));
    InMux I__5331 (
            .O(N__24168),
            .I(N__24150));
    InMux I__5330 (
            .O(N__24165),
            .I(N__24150));
    Span4Mux_h I__5329 (
            .O(N__24162),
            .I(N__24145));
    LocalMux I__5328 (
            .O(N__24159),
            .I(N__24145));
    InMux I__5327 (
            .O(N__24158),
            .I(N__24140));
    InMux I__5326 (
            .O(N__24157),
            .I(N__24140));
    LocalMux I__5325 (
            .O(N__24150),
            .I(\Lab_UT.dictrl.un2_dicAlarmTrig ));
    Odrv4 I__5324 (
            .O(N__24145),
            .I(\Lab_UT.dictrl.un2_dicAlarmTrig ));
    LocalMux I__5323 (
            .O(N__24140),
            .I(\Lab_UT.dictrl.un2_dicAlarmTrig ));
    InMux I__5322 (
            .O(N__24133),
            .I(N__24130));
    LocalMux I__5321 (
            .O(N__24130),
            .I(\Lab_UT.dictrl.N_186 ));
    CascadeMux I__5320 (
            .O(N__24127),
            .I(N__24123));
    InMux I__5319 (
            .O(N__24126),
            .I(N__24113));
    InMux I__5318 (
            .O(N__24123),
            .I(N__24113));
    InMux I__5317 (
            .O(N__24122),
            .I(N__24113));
    CascadeMux I__5316 (
            .O(N__24121),
            .I(N__24110));
    CascadeMux I__5315 (
            .O(N__24120),
            .I(N__24107));
    LocalMux I__5314 (
            .O(N__24113),
            .I(N__24104));
    InMux I__5313 (
            .O(N__24110),
            .I(N__24101));
    InMux I__5312 (
            .O(N__24107),
            .I(N__24098));
    Span4Mux_h I__5311 (
            .O(N__24104),
            .I(N__24095));
    LocalMux I__5310 (
            .O(N__24101),
            .I(\Lab_UT.dictrl.nextState_al_0_0 ));
    LocalMux I__5309 (
            .O(N__24098),
            .I(\Lab_UT.dictrl.nextState_al_0_0 ));
    Odrv4 I__5308 (
            .O(N__24095),
            .I(\Lab_UT.dictrl.nextState_al_0_0 ));
    CascadeMux I__5307 (
            .O(N__24088),
            .I(\Lab_UT.dictrl.N_186_cascade_ ));
    InMux I__5306 (
            .O(N__24085),
            .I(N__24081));
    InMux I__5305 (
            .O(N__24084),
            .I(N__24078));
    LocalMux I__5304 (
            .O(N__24081),
            .I(\Lab_UT.dictrl.nextState_al_1_0_0_1 ));
    LocalMux I__5303 (
            .O(N__24078),
            .I(\Lab_UT.dictrl.nextState_al_1_0_0_1 ));
    CascadeMux I__5302 (
            .O(N__24073),
            .I(N__24069));
    InMux I__5301 (
            .O(N__24072),
            .I(N__24061));
    InMux I__5300 (
            .O(N__24069),
            .I(N__24061));
    InMux I__5299 (
            .O(N__24068),
            .I(N__24061));
    LocalMux I__5298 (
            .O(N__24061),
            .I(\Lab_UT.dictrl.currState_alZ0Z_0 ));
    InMux I__5297 (
            .O(N__24058),
            .I(N__24047));
    InMux I__5296 (
            .O(N__24057),
            .I(N__24047));
    InMux I__5295 (
            .O(N__24056),
            .I(N__24044));
    InMux I__5294 (
            .O(N__24055),
            .I(N__24035));
    InMux I__5293 (
            .O(N__24054),
            .I(N__24035));
    InMux I__5292 (
            .O(N__24053),
            .I(N__24035));
    InMux I__5291 (
            .O(N__24052),
            .I(N__24035));
    LocalMux I__5290 (
            .O(N__24047),
            .I(\Lab_UT.dictrl.currState_alZ0Z_1 ));
    LocalMux I__5289 (
            .O(N__24044),
            .I(\Lab_UT.dictrl.currState_alZ0Z_1 ));
    LocalMux I__5288 (
            .O(N__24035),
            .I(\Lab_UT.dictrl.currState_alZ0Z_1 ));
    CascadeMux I__5287 (
            .O(N__24028),
            .I(N__24025));
    InMux I__5286 (
            .O(N__24025),
            .I(N__24022));
    LocalMux I__5285 (
            .O(N__24022),
            .I(N__24019));
    Span12Mux_s11_h I__5284 (
            .O(N__24019),
            .I(N__24016));
    Odrv12 I__5283 (
            .O(N__24016),
            .I(\Lab_UT.dictrl.currState_i_5_1 ));
    InMux I__5282 (
            .O(N__24013),
            .I(N__24008));
    CascadeMux I__5281 (
            .O(N__24012),
            .I(N__24000));
    InMux I__5280 (
            .O(N__24011),
            .I(N__23997));
    LocalMux I__5279 (
            .O(N__24008),
            .I(N__23994));
    InMux I__5278 (
            .O(N__24007),
            .I(N__23991));
    InMux I__5277 (
            .O(N__24006),
            .I(N__23988));
    InMux I__5276 (
            .O(N__24005),
            .I(N__23985));
    InMux I__5275 (
            .O(N__24004),
            .I(N__23982));
    InMux I__5274 (
            .O(N__24003),
            .I(N__23977));
    InMux I__5273 (
            .O(N__24000),
            .I(N__23977));
    LocalMux I__5272 (
            .O(N__23997),
            .I(N__23973));
    Span4Mux_v I__5271 (
            .O(N__23994),
            .I(N__23969));
    LocalMux I__5270 (
            .O(N__23991),
            .I(N__23966));
    LocalMux I__5269 (
            .O(N__23988),
            .I(N__23963));
    LocalMux I__5268 (
            .O(N__23985),
            .I(N__23960));
    LocalMux I__5267 (
            .O(N__23982),
            .I(N__23955));
    LocalMux I__5266 (
            .O(N__23977),
            .I(N__23955));
    InMux I__5265 (
            .O(N__23976),
            .I(N__23952));
    Span4Mux_v I__5264 (
            .O(N__23973),
            .I(N__23949));
    InMux I__5263 (
            .O(N__23972),
            .I(N__23946));
    Span4Mux_h I__5262 (
            .O(N__23969),
            .I(N__23937));
    Span4Mux_v I__5261 (
            .O(N__23966),
            .I(N__23937));
    Span4Mux_v I__5260 (
            .O(N__23963),
            .I(N__23937));
    Span4Mux_v I__5259 (
            .O(N__23960),
            .I(N__23937));
    Span4Mux_v I__5258 (
            .O(N__23955),
            .I(N__23934));
    LocalMux I__5257 (
            .O(N__23952),
            .I(\Lab_UT.dictrl.currState_i_5_0 ));
    Odrv4 I__5256 (
            .O(N__23949),
            .I(\Lab_UT.dictrl.currState_i_5_0 ));
    LocalMux I__5255 (
            .O(N__23946),
            .I(\Lab_UT.dictrl.currState_i_5_0 ));
    Odrv4 I__5254 (
            .O(N__23937),
            .I(\Lab_UT.dictrl.currState_i_5_0 ));
    Odrv4 I__5253 (
            .O(N__23934),
            .I(\Lab_UT.dictrl.currState_i_5_0 ));
    CascadeMux I__5252 (
            .O(N__23923),
            .I(\Lab_UT.dictrl.un1_currState_8_u_ns_1_cascade_ ));
    SRMux I__5251 (
            .O(N__23920),
            .I(N__23917));
    LocalMux I__5250 (
            .O(N__23917),
            .I(N__23914));
    Sp12to4 I__5249 (
            .O(N__23914),
            .I(N__23910));
    InMux I__5248 (
            .O(N__23913),
            .I(N__23907));
    Odrv12 I__5247 (
            .O(N__23910),
            .I(\Lab_UT.dictrl.currState_ret_7_RNI03VHZ0Z1 ));
    LocalMux I__5246 (
            .O(N__23907),
            .I(\Lab_UT.dictrl.currState_ret_7_RNI03VHZ0Z1 ));
    CascadeMux I__5245 (
            .O(N__23902),
            .I(\Lab_UT.dictrl.un1_currState_inv_1_cascade_ ));
    SRMux I__5244 (
            .O(N__23899),
            .I(N__23895));
    InMux I__5243 (
            .O(N__23898),
            .I(N__23892));
    LocalMux I__5242 (
            .O(N__23895),
            .I(N__23889));
    LocalMux I__5241 (
            .O(N__23892),
            .I(N__23886));
    Span4Mux_h I__5240 (
            .O(N__23889),
            .I(N__23883));
    Span4Mux_v I__5239 (
            .O(N__23886),
            .I(N__23880));
    Span4Mux_v I__5238 (
            .O(N__23883),
            .I(N__23877));
    Span4Mux_h I__5237 (
            .O(N__23880),
            .I(N__23874));
    Odrv4 I__5236 (
            .O(N__23877),
            .I(\Lab_UT.dictrl.currState_0_ret_1_RNIPH7FZ0Z1 ));
    Odrv4 I__5235 (
            .O(N__23874),
            .I(\Lab_UT.dictrl.currState_0_ret_1_RNIPH7FZ0Z1 ));
    InMux I__5234 (
            .O(N__23869),
            .I(N__23866));
    LocalMux I__5233 (
            .O(N__23866),
            .I(N__23863));
    Odrv12 I__5232 (
            .O(N__23863),
            .I(\Lab_UT.dictrl.r_dicLdMtens14_1 ));
    InMux I__5231 (
            .O(N__23860),
            .I(N__23857));
    LocalMux I__5230 (
            .O(N__23857),
            .I(N__23851));
    InMux I__5229 (
            .O(N__23856),
            .I(N__23846));
    InMux I__5228 (
            .O(N__23855),
            .I(N__23846));
    InMux I__5227 (
            .O(N__23854),
            .I(N__23843));
    Span4Mux_h I__5226 (
            .O(N__23851),
            .I(N__23836));
    LocalMux I__5225 (
            .O(N__23846),
            .I(N__23836));
    LocalMux I__5224 (
            .O(N__23843),
            .I(N__23836));
    Odrv4 I__5223 (
            .O(N__23836),
            .I(\Lab_UT.dictrl.r_Sone_init5_1 ));
    CascadeMux I__5222 (
            .O(N__23833),
            .I(N__23828));
    InMux I__5221 (
            .O(N__23832),
            .I(N__23819));
    InMux I__5220 (
            .O(N__23831),
            .I(N__23819));
    InMux I__5219 (
            .O(N__23828),
            .I(N__23807));
    InMux I__5218 (
            .O(N__23827),
            .I(N__23807));
    InMux I__5217 (
            .O(N__23826),
            .I(N__23804));
    InMux I__5216 (
            .O(N__23825),
            .I(N__23799));
    InMux I__5215 (
            .O(N__23824),
            .I(N__23799));
    LocalMux I__5214 (
            .O(N__23819),
            .I(N__23795));
    InMux I__5213 (
            .O(N__23818),
            .I(N__23792));
    InMux I__5212 (
            .O(N__23817),
            .I(N__23789));
    InMux I__5211 (
            .O(N__23816),
            .I(N__23786));
    InMux I__5210 (
            .O(N__23815),
            .I(N__23781));
    InMux I__5209 (
            .O(N__23814),
            .I(N__23778));
    InMux I__5208 (
            .O(N__23813),
            .I(N__23772));
    InMux I__5207 (
            .O(N__23812),
            .I(N__23769));
    LocalMux I__5206 (
            .O(N__23807),
            .I(N__23764));
    LocalMux I__5205 (
            .O(N__23804),
            .I(N__23764));
    LocalMux I__5204 (
            .O(N__23799),
            .I(N__23761));
    InMux I__5203 (
            .O(N__23798),
            .I(N__23758));
    Span4Mux_v I__5202 (
            .O(N__23795),
            .I(N__23749));
    LocalMux I__5201 (
            .O(N__23792),
            .I(N__23749));
    LocalMux I__5200 (
            .O(N__23789),
            .I(N__23749));
    LocalMux I__5199 (
            .O(N__23786),
            .I(N__23749));
    InMux I__5198 (
            .O(N__23785),
            .I(N__23744));
    InMux I__5197 (
            .O(N__23784),
            .I(N__23744));
    LocalMux I__5196 (
            .O(N__23781),
            .I(N__23741));
    LocalMux I__5195 (
            .O(N__23778),
            .I(N__23738));
    InMux I__5194 (
            .O(N__23777),
            .I(N__23731));
    InMux I__5193 (
            .O(N__23776),
            .I(N__23731));
    InMux I__5192 (
            .O(N__23775),
            .I(N__23731));
    LocalMux I__5191 (
            .O(N__23772),
            .I(N__23724));
    LocalMux I__5190 (
            .O(N__23769),
            .I(N__23724));
    Span4Mux_h I__5189 (
            .O(N__23764),
            .I(N__23724));
    Span4Mux_v I__5188 (
            .O(N__23761),
            .I(N__23721));
    LocalMux I__5187 (
            .O(N__23758),
            .I(N__23716));
    Span4Mux_h I__5186 (
            .O(N__23749),
            .I(N__23716));
    LocalMux I__5185 (
            .O(N__23744),
            .I(N__23709));
    Span4Mux_v I__5184 (
            .O(N__23741),
            .I(N__23709));
    Span4Mux_s3_h I__5183 (
            .O(N__23738),
            .I(N__23709));
    LocalMux I__5182 (
            .O(N__23731),
            .I(N__23704));
    Span4Mux_h I__5181 (
            .O(N__23724),
            .I(N__23704));
    Span4Mux_h I__5180 (
            .O(N__23721),
            .I(N__23699));
    Span4Mux_v I__5179 (
            .O(N__23716),
            .I(N__23699));
    Span4Mux_h I__5178 (
            .O(N__23709),
            .I(N__23696));
    Span4Mux_v I__5177 (
            .O(N__23704),
            .I(N__23693));
    Odrv4 I__5176 (
            .O(N__23699),
            .I(\Lab_UT.dictrl.currStateZ0Z_3 ));
    Odrv4 I__5175 (
            .O(N__23696),
            .I(\Lab_UT.dictrl.currStateZ0Z_3 ));
    Odrv4 I__5174 (
            .O(N__23693),
            .I(\Lab_UT.dictrl.currStateZ0Z_3 ));
    InMux I__5173 (
            .O(N__23686),
            .I(N__23682));
    InMux I__5172 (
            .O(N__23685),
            .I(N__23679));
    LocalMux I__5171 (
            .O(N__23682),
            .I(\Lab_UT.dictrl.un1_currState_inv_1 ));
    LocalMux I__5170 (
            .O(N__23679),
            .I(\Lab_UT.dictrl.un1_currState_inv_1 ));
    CascadeMux I__5169 (
            .O(N__23674),
            .I(\Lab_UT.dictrl.N_201_cascade_ ));
    SRMux I__5168 (
            .O(N__23671),
            .I(N__23665));
    InMux I__5167 (
            .O(N__23670),
            .I(N__23665));
    LocalMux I__5166 (
            .O(N__23665),
            .I(N__23662));
    Span4Mux_h I__5165 (
            .O(N__23662),
            .I(N__23659));
    Odrv4 I__5164 (
            .O(N__23659),
            .I(\Lab_UT.dictrl.currState_2_RNIOB6H1Z0Z_2 ));
    InMux I__5163 (
            .O(N__23656),
            .I(N__23647));
    InMux I__5162 (
            .O(N__23655),
            .I(N__23647));
    InMux I__5161 (
            .O(N__23654),
            .I(N__23647));
    LocalMux I__5160 (
            .O(N__23647),
            .I(N__23642));
    InMux I__5159 (
            .O(N__23646),
            .I(N__23639));
    InMux I__5158 (
            .O(N__23645),
            .I(N__23634));
    Span4Mux_h I__5157 (
            .O(N__23642),
            .I(N__23631));
    LocalMux I__5156 (
            .O(N__23639),
            .I(N__23628));
    InMux I__5155 (
            .O(N__23638),
            .I(N__23623));
    InMux I__5154 (
            .O(N__23637),
            .I(N__23623));
    LocalMux I__5153 (
            .O(N__23634),
            .I(\Lab_UT.dictrl.r_dicAlarmTrigZ0 ));
    Odrv4 I__5152 (
            .O(N__23631),
            .I(\Lab_UT.dictrl.r_dicAlarmTrigZ0 ));
    Odrv4 I__5151 (
            .O(N__23628),
            .I(\Lab_UT.dictrl.r_dicAlarmTrigZ0 ));
    LocalMux I__5150 (
            .O(N__23623),
            .I(\Lab_UT.dictrl.r_dicAlarmTrigZ0 ));
    InMux I__5149 (
            .O(N__23614),
            .I(N__23611));
    LocalMux I__5148 (
            .O(N__23611),
            .I(N__23608));
    Odrv12 I__5147 (
            .O(N__23608),
            .I(\Lab_UT.displayAlarmZ0Z_5 ));
    InMux I__5146 (
            .O(N__23605),
            .I(N__23602));
    LocalMux I__5145 (
            .O(N__23602),
            .I(\Lab_UT.dictrl.nextState_al_1 ));
    CascadeMux I__5144 (
            .O(N__23599),
            .I(\Lab_UT.dictrl.nextState_al_1_cascade_ ));
    CascadeMux I__5143 (
            .O(N__23596),
            .I(N__23592));
    InMux I__5142 (
            .O(N__23595),
            .I(N__23589));
    InMux I__5141 (
            .O(N__23592),
            .I(N__23586));
    LocalMux I__5140 (
            .O(N__23589),
            .I(\Lab_UT.dictrl.un2_dicAlarmTrig_i_6 ));
    LocalMux I__5139 (
            .O(N__23586),
            .I(\Lab_UT.dictrl.un2_dicAlarmTrig_i_6 ));
    InMux I__5138 (
            .O(N__23581),
            .I(N__23578));
    LocalMux I__5137 (
            .O(N__23578),
            .I(\Lab_UT.dictrl.nextState_al_latmux_1 ));
    CascadeMux I__5136 (
            .O(N__23575),
            .I(\Lab_UT.dictrl.nextState_al_latmux_1_cascade_ ));
    InMux I__5135 (
            .O(N__23572),
            .I(N__23566));
    InMux I__5134 (
            .O(N__23571),
            .I(N__23566));
    LocalMux I__5133 (
            .O(N__23566),
            .I(\Lab_UT.dictrl.nextState_alZ0Z_0 ));
    InMux I__5132 (
            .O(N__23563),
            .I(N__23560));
    LocalMux I__5131 (
            .O(N__23560),
            .I(\Lab_UT.didp.Stens_subtractor.un1_q_axb0 ));
    InMux I__5130 (
            .O(N__23557),
            .I(N__23554));
    LocalMux I__5129 (
            .O(N__23554),
            .I(\Lab_UT.didp.Stens_subtractor.q_RNO_0_0_3 ));
    InMux I__5128 (
            .O(N__23551),
            .I(N__23542));
    InMux I__5127 (
            .O(N__23550),
            .I(N__23542));
    InMux I__5126 (
            .O(N__23549),
            .I(N__23542));
    LocalMux I__5125 (
            .O(N__23542),
            .I(\Lab_UT.didp.Stens_subtractor.N_86 ));
    InMux I__5124 (
            .O(N__23539),
            .I(N__23536));
    LocalMux I__5123 (
            .O(N__23536),
            .I(\Lab_UT.didp.Stens_subtractor.q_RNO_0_1_2 ));
    CascadeMux I__5122 (
            .O(N__23533),
            .I(\Lab_UT.didp.q_RNIDDF11_3_cascade_ ));
    IoInMux I__5121 (
            .O(N__23530),
            .I(N__23527));
    LocalMux I__5120 (
            .O(N__23527),
            .I(N__23524));
    Span4Mux_s3_h I__5119 (
            .O(N__23524),
            .I(N__23521));
    Odrv4 I__5118 (
            .O(N__23521),
            .I(led_c_3));
    InMux I__5117 (
            .O(N__23518),
            .I(N__23515));
    LocalMux I__5116 (
            .O(N__23515),
            .I(\Lab_UT.didp.q_RNI1TVP_3 ));
    InMux I__5115 (
            .O(N__23512),
            .I(N__23509));
    LocalMux I__5114 (
            .O(N__23509),
            .I(\Lab_UT.didp.q_RNIBBF11_2 ));
    InMux I__5113 (
            .O(N__23506),
            .I(N__23503));
    LocalMux I__5112 (
            .O(N__23503),
            .I(N__23500));
    Span4Mux_h I__5111 (
            .O(N__23500),
            .I(N__23497));
    Odrv4 I__5110 (
            .O(N__23497),
            .I(\Lab_UT.didp.q_RNIVQVP_2 ));
    IoInMux I__5109 (
            .O(N__23494),
            .I(N__23491));
    LocalMux I__5108 (
            .O(N__23491),
            .I(N__23488));
    Span4Mux_s2_h I__5107 (
            .O(N__23488),
            .I(N__23485));
    Odrv4 I__5106 (
            .O(N__23485),
            .I(led_c_2));
    InMux I__5105 (
            .O(N__23482),
            .I(N__23479));
    LocalMux I__5104 (
            .O(N__23479),
            .I(N__23473));
    InMux I__5103 (
            .O(N__23478),
            .I(N__23470));
    InMux I__5102 (
            .O(N__23477),
            .I(N__23465));
    InMux I__5101 (
            .O(N__23476),
            .I(N__23465));
    Odrv4 I__5100 (
            .O(N__23473),
            .I(\Lab_UT.dictrl.r_Sone_init5 ));
    LocalMux I__5099 (
            .O(N__23470),
            .I(\Lab_UT.dictrl.r_Sone_init5 ));
    LocalMux I__5098 (
            .O(N__23465),
            .I(\Lab_UT.dictrl.r_Sone_init5 ));
    CascadeMux I__5097 (
            .O(N__23458),
            .I(N__23449));
    CascadeMux I__5096 (
            .O(N__23457),
            .I(N__23441));
    InMux I__5095 (
            .O(N__23456),
            .I(N__23432));
    InMux I__5094 (
            .O(N__23455),
            .I(N__23423));
    InMux I__5093 (
            .O(N__23454),
            .I(N__23423));
    InMux I__5092 (
            .O(N__23453),
            .I(N__23423));
    InMux I__5091 (
            .O(N__23452),
            .I(N__23415));
    InMux I__5090 (
            .O(N__23449),
            .I(N__23415));
    InMux I__5089 (
            .O(N__23448),
            .I(N__23415));
    InMux I__5088 (
            .O(N__23447),
            .I(N__23412));
    InMux I__5087 (
            .O(N__23446),
            .I(N__23405));
    InMux I__5086 (
            .O(N__23445),
            .I(N__23405));
    InMux I__5085 (
            .O(N__23444),
            .I(N__23405));
    InMux I__5084 (
            .O(N__23441),
            .I(N__23402));
    InMux I__5083 (
            .O(N__23440),
            .I(N__23397));
    InMux I__5082 (
            .O(N__23439),
            .I(N__23397));
    InMux I__5081 (
            .O(N__23438),
            .I(N__23390));
    InMux I__5080 (
            .O(N__23437),
            .I(N__23390));
    InMux I__5079 (
            .O(N__23436),
            .I(N__23390));
    InMux I__5078 (
            .O(N__23435),
            .I(N__23385));
    LocalMux I__5077 (
            .O(N__23432),
            .I(N__23382));
    InMux I__5076 (
            .O(N__23431),
            .I(N__23378));
    InMux I__5075 (
            .O(N__23430),
            .I(N__23372));
    LocalMux I__5074 (
            .O(N__23423),
            .I(N__23369));
    InMux I__5073 (
            .O(N__23422),
            .I(N__23366));
    LocalMux I__5072 (
            .O(N__23415),
            .I(N__23363));
    LocalMux I__5071 (
            .O(N__23412),
            .I(N__23358));
    LocalMux I__5070 (
            .O(N__23405),
            .I(N__23358));
    LocalMux I__5069 (
            .O(N__23402),
            .I(N__23351));
    LocalMux I__5068 (
            .O(N__23397),
            .I(N__23351));
    LocalMux I__5067 (
            .O(N__23390),
            .I(N__23351));
    InMux I__5066 (
            .O(N__23389),
            .I(N__23346));
    InMux I__5065 (
            .O(N__23388),
            .I(N__23346));
    LocalMux I__5064 (
            .O(N__23385),
            .I(N__23337));
    Span4Mux_s3_h I__5063 (
            .O(N__23382),
            .I(N__23334));
    InMux I__5062 (
            .O(N__23381),
            .I(N__23331));
    LocalMux I__5061 (
            .O(N__23378),
            .I(N__23328));
    InMux I__5060 (
            .O(N__23377),
            .I(N__23321));
    InMux I__5059 (
            .O(N__23376),
            .I(N__23321));
    InMux I__5058 (
            .O(N__23375),
            .I(N__23318));
    LocalMux I__5057 (
            .O(N__23372),
            .I(N__23315));
    Span4Mux_v I__5056 (
            .O(N__23369),
            .I(N__23308));
    LocalMux I__5055 (
            .O(N__23366),
            .I(N__23308));
    Span4Mux_h I__5054 (
            .O(N__23363),
            .I(N__23308));
    Span4Mux_v I__5053 (
            .O(N__23358),
            .I(N__23301));
    Span4Mux_h I__5052 (
            .O(N__23351),
            .I(N__23301));
    LocalMux I__5051 (
            .O(N__23346),
            .I(N__23301));
    InMux I__5050 (
            .O(N__23345),
            .I(N__23298));
    InMux I__5049 (
            .O(N__23344),
            .I(N__23295));
    InMux I__5048 (
            .O(N__23343),
            .I(N__23286));
    InMux I__5047 (
            .O(N__23342),
            .I(N__23286));
    InMux I__5046 (
            .O(N__23341),
            .I(N__23286));
    InMux I__5045 (
            .O(N__23340),
            .I(N__23286));
    Span4Mux_h I__5044 (
            .O(N__23337),
            .I(N__23277));
    Span4Mux_h I__5043 (
            .O(N__23334),
            .I(N__23277));
    LocalMux I__5042 (
            .O(N__23331),
            .I(N__23277));
    Span4Mux_v I__5041 (
            .O(N__23328),
            .I(N__23277));
    InMux I__5040 (
            .O(N__23327),
            .I(N__23272));
    InMux I__5039 (
            .O(N__23326),
            .I(N__23272));
    LocalMux I__5038 (
            .O(N__23321),
            .I(N__23261));
    LocalMux I__5037 (
            .O(N__23318),
            .I(N__23261));
    Span4Mux_h I__5036 (
            .O(N__23315),
            .I(N__23261));
    Span4Mux_h I__5035 (
            .O(N__23308),
            .I(N__23261));
    Span4Mux_h I__5034 (
            .O(N__23301),
            .I(N__23261));
    LocalMux I__5033 (
            .O(N__23298),
            .I(Lab_UT_dictrl_r_Sone_init17));
    LocalMux I__5032 (
            .O(N__23295),
            .I(Lab_UT_dictrl_r_Sone_init17));
    LocalMux I__5031 (
            .O(N__23286),
            .I(Lab_UT_dictrl_r_Sone_init17));
    Odrv4 I__5030 (
            .O(N__23277),
            .I(Lab_UT_dictrl_r_Sone_init17));
    LocalMux I__5029 (
            .O(N__23272),
            .I(Lab_UT_dictrl_r_Sone_init17));
    Odrv4 I__5028 (
            .O(N__23261),
            .I(Lab_UT_dictrl_r_Sone_init17));
    InMux I__5027 (
            .O(N__23248),
            .I(N__23241));
    InMux I__5026 (
            .O(N__23247),
            .I(N__23241));
    InMux I__5025 (
            .O(N__23246),
            .I(N__23236));
    LocalMux I__5024 (
            .O(N__23241),
            .I(N__23229));
    InMux I__5023 (
            .O(N__23240),
            .I(N__23224));
    InMux I__5022 (
            .O(N__23239),
            .I(N__23224));
    LocalMux I__5021 (
            .O(N__23236),
            .I(N__23217));
    InMux I__5020 (
            .O(N__23235),
            .I(N__23214));
    InMux I__5019 (
            .O(N__23234),
            .I(N__23207));
    InMux I__5018 (
            .O(N__23233),
            .I(N__23207));
    InMux I__5017 (
            .O(N__23232),
            .I(N__23207));
    Span4Mux_s1_v I__5016 (
            .O(N__23229),
            .I(N__23202));
    LocalMux I__5015 (
            .O(N__23224),
            .I(N__23202));
    InMux I__5014 (
            .O(N__23223),
            .I(N__23199));
    InMux I__5013 (
            .O(N__23222),
            .I(N__23192));
    InMux I__5012 (
            .O(N__23221),
            .I(N__23192));
    InMux I__5011 (
            .O(N__23220),
            .I(N__23192));
    Span4Mux_v I__5010 (
            .O(N__23217),
            .I(N__23187));
    LocalMux I__5009 (
            .O(N__23214),
            .I(N__23187));
    LocalMux I__5008 (
            .O(N__23207),
            .I(\Lab_UT.uu0.un4_l_count_0 ));
    Odrv4 I__5007 (
            .O(N__23202),
            .I(\Lab_UT.uu0.un4_l_count_0 ));
    LocalMux I__5006 (
            .O(N__23199),
            .I(\Lab_UT.uu0.un4_l_count_0 ));
    LocalMux I__5005 (
            .O(N__23192),
            .I(\Lab_UT.uu0.un4_l_count_0 ));
    Odrv4 I__5004 (
            .O(N__23187),
            .I(\Lab_UT.uu0.un4_l_count_0 ));
    CascadeMux I__5003 (
            .O(N__23176),
            .I(N__23171));
    InMux I__5002 (
            .O(N__23175),
            .I(N__23163));
    InMux I__5001 (
            .O(N__23174),
            .I(N__23163));
    InMux I__5000 (
            .O(N__23171),
            .I(N__23163));
    CascadeMux I__4999 (
            .O(N__23170),
            .I(N__23158));
    LocalMux I__4998 (
            .O(N__23163),
            .I(N__23154));
    InMux I__4997 (
            .O(N__23162),
            .I(N__23147));
    InMux I__4996 (
            .O(N__23161),
            .I(N__23147));
    InMux I__4995 (
            .O(N__23158),
            .I(N__23147));
    InMux I__4994 (
            .O(N__23157),
            .I(N__23144));
    Span4Mux_h I__4993 (
            .O(N__23154),
            .I(N__23141));
    LocalMux I__4992 (
            .O(N__23147),
            .I(N__23138));
    LocalMux I__4991 (
            .O(N__23144),
            .I(\Lab_UT.halfPulse ));
    Odrv4 I__4990 (
            .O(N__23141),
            .I(\Lab_UT.halfPulse ));
    Odrv4 I__4989 (
            .O(N__23138),
            .I(\Lab_UT.halfPulse ));
    InMux I__4988 (
            .O(N__23131),
            .I(N__23127));
    InMux I__4987 (
            .O(N__23130),
            .I(N__23124));
    LocalMux I__4986 (
            .O(N__23127),
            .I(N__23121));
    LocalMux I__4985 (
            .O(N__23124),
            .I(N__23118));
    Odrv12 I__4984 (
            .O(N__23121),
            .I(\Lab_UT.displayAlarmZ0Z_1 ));
    Odrv4 I__4983 (
            .O(N__23118),
            .I(\Lab_UT.displayAlarmZ0Z_1 ));
    CascadeMux I__4982 (
            .O(N__23113),
            .I(N__23109));
    CascadeMux I__4981 (
            .O(N__23112),
            .I(N__23106));
    InMux I__4980 (
            .O(N__23109),
            .I(N__23102));
    InMux I__4979 (
            .O(N__23106),
            .I(N__23097));
    InMux I__4978 (
            .O(N__23105),
            .I(N__23097));
    LocalMux I__4977 (
            .O(N__23102),
            .I(\Lab_UT.dicLdStens ));
    LocalMux I__4976 (
            .O(N__23097),
            .I(\Lab_UT.dicLdStens ));
    InMux I__4975 (
            .O(N__23092),
            .I(N__23087));
    InMux I__4974 (
            .O(N__23091),
            .I(N__23082));
    InMux I__4973 (
            .O(N__23090),
            .I(N__23082));
    LocalMux I__4972 (
            .O(N__23087),
            .I(\Lab_UT.dicLdStens_latmux ));
    LocalMux I__4971 (
            .O(N__23082),
            .I(\Lab_UT.dicLdStens_latmux ));
    InMux I__4970 (
            .O(N__23077),
            .I(N__23072));
    InMux I__4969 (
            .O(N__23076),
            .I(N__23069));
    InMux I__4968 (
            .O(N__23075),
            .I(N__23066));
    LocalMux I__4967 (
            .O(N__23072),
            .I(\Lab_UT.di_ASones_0 ));
    LocalMux I__4966 (
            .O(N__23069),
            .I(\Lab_UT.di_ASones_0 ));
    LocalMux I__4965 (
            .O(N__23066),
            .I(\Lab_UT.di_ASones_0 ));
    InMux I__4964 (
            .O(N__23059),
            .I(N__23054));
    InMux I__4963 (
            .O(N__23058),
            .I(N__23051));
    InMux I__4962 (
            .O(N__23057),
            .I(N__23048));
    LocalMux I__4961 (
            .O(N__23054),
            .I(N__23045));
    LocalMux I__4960 (
            .O(N__23051),
            .I(\Lab_UT.di_ASones_1 ));
    LocalMux I__4959 (
            .O(N__23048),
            .I(\Lab_UT.di_ASones_1 ));
    Odrv4 I__4958 (
            .O(N__23045),
            .I(\Lab_UT.di_ASones_1 ));
    InMux I__4957 (
            .O(N__23038),
            .I(N__23033));
    InMux I__4956 (
            .O(N__23037),
            .I(N__23030));
    InMux I__4955 (
            .O(N__23036),
            .I(N__23027));
    LocalMux I__4954 (
            .O(N__23033),
            .I(\Lab_UT.di_ASones_2 ));
    LocalMux I__4953 (
            .O(N__23030),
            .I(\Lab_UT.di_ASones_2 ));
    LocalMux I__4952 (
            .O(N__23027),
            .I(\Lab_UT.di_ASones_2 ));
    CascadeMux I__4951 (
            .O(N__23020),
            .I(N__23015));
    InMux I__4950 (
            .O(N__23019),
            .I(N__23011));
    InMux I__4949 (
            .O(N__23018),
            .I(N__23008));
    InMux I__4948 (
            .O(N__23015),
            .I(N__23003));
    InMux I__4947 (
            .O(N__23014),
            .I(N__23003));
    LocalMux I__4946 (
            .O(N__23011),
            .I(N__22998));
    LocalMux I__4945 (
            .O(N__23008),
            .I(N__22998));
    LocalMux I__4944 (
            .O(N__23003),
            .I(N__22995));
    Span4Mux_h I__4943 (
            .O(N__22998),
            .I(N__22992));
    Span4Mux_h I__4942 (
            .O(N__22995),
            .I(N__22989));
    Odrv4 I__4941 (
            .O(N__22992),
            .I(\Lab_UT.ld_enable_AMtens ));
    Odrv4 I__4940 (
            .O(N__22989),
            .I(\Lab_UT.ld_enable_AMtens ));
    InMux I__4939 (
            .O(N__22984),
            .I(N__22980));
    InMux I__4938 (
            .O(N__22983),
            .I(N__22976));
    LocalMux I__4937 (
            .O(N__22980),
            .I(N__22973));
    InMux I__4936 (
            .O(N__22979),
            .I(N__22970));
    LocalMux I__4935 (
            .O(N__22976),
            .I(\Lab_UT.di_AStens_3 ));
    Odrv4 I__4934 (
            .O(N__22973),
            .I(\Lab_UT.di_AStens_3 ));
    LocalMux I__4933 (
            .O(N__22970),
            .I(\Lab_UT.di_AStens_3 ));
    InMux I__4932 (
            .O(N__22963),
            .I(N__22954));
    InMux I__4931 (
            .O(N__22962),
            .I(N__22954));
    InMux I__4930 (
            .O(N__22961),
            .I(N__22954));
    LocalMux I__4929 (
            .O(N__22954),
            .I(N__22950));
    InMux I__4928 (
            .O(N__22953),
            .I(N__22947));
    Span4Mux_v I__4927 (
            .O(N__22950),
            .I(N__22944));
    LocalMux I__4926 (
            .O(N__22947),
            .I(N__22941));
    Span4Mux_v I__4925 (
            .O(N__22944),
            .I(N__22938));
    Span4Mux_h I__4924 (
            .O(N__22941),
            .I(N__22935));
    Odrv4 I__4923 (
            .O(N__22938),
            .I(\Lab_UT.ld_enable_ASones ));
    Odrv4 I__4922 (
            .O(N__22935),
            .I(\Lab_UT.ld_enable_ASones ));
    InMux I__4921 (
            .O(N__22930),
            .I(N__22926));
    InMux I__4920 (
            .O(N__22929),
            .I(N__22922));
    LocalMux I__4919 (
            .O(N__22926),
            .I(N__22919));
    InMux I__4918 (
            .O(N__22925),
            .I(N__22916));
    LocalMux I__4917 (
            .O(N__22922),
            .I(\Lab_UT.di_ASones_3 ));
    Odrv4 I__4916 (
            .O(N__22919),
            .I(\Lab_UT.di_ASones_3 ));
    LocalMux I__4915 (
            .O(N__22916),
            .I(\Lab_UT.di_ASones_3 ));
    InMux I__4914 (
            .O(N__22909),
            .I(N__22897));
    InMux I__4913 (
            .O(N__22908),
            .I(N__22897));
    InMux I__4912 (
            .O(N__22907),
            .I(N__22897));
    InMux I__4911 (
            .O(N__22906),
            .I(N__22897));
    LocalMux I__4910 (
            .O(N__22897),
            .I(N__22894));
    Span4Mux_v I__4909 (
            .O(N__22894),
            .I(N__22891));
    Odrv4 I__4908 (
            .O(N__22891),
            .I(\Lab_UT.ld_enable_AStens ));
    InMux I__4907 (
            .O(N__22888),
            .I(N__22885));
    LocalMux I__4906 (
            .O(N__22885),
            .I(\Lab_UT.display.dOutP_0_iv_i_1_1 ));
    CascadeMux I__4905 (
            .O(N__22882),
            .I(N__22878));
    CascadeMux I__4904 (
            .O(N__22881),
            .I(N__22875));
    InMux I__4903 (
            .O(N__22878),
            .I(N__22864));
    InMux I__4902 (
            .O(N__22875),
            .I(N__22864));
    InMux I__4901 (
            .O(N__22874),
            .I(N__22864));
    InMux I__4900 (
            .O(N__22873),
            .I(N__22864));
    LocalMux I__4899 (
            .O(N__22864),
            .I(\Lab_UT.display.N_150 ));
    CascadeMux I__4898 (
            .O(N__22861),
            .I(\Lab_UT.display.N_101_cascade_ ));
    InMux I__4897 (
            .O(N__22858),
            .I(N__22855));
    LocalMux I__4896 (
            .O(N__22855),
            .I(N__22851));
    InMux I__4895 (
            .O(N__22854),
            .I(N__22848));
    Odrv4 I__4894 (
            .O(N__22851),
            .I(\Lab_UT.display.N_88 ));
    LocalMux I__4893 (
            .O(N__22848),
            .I(\Lab_UT.display.N_88 ));
    CascadeMux I__4892 (
            .O(N__22843),
            .I(\Lab_UT.display.dOutP_0_iv_i_0_3_cascade_ ));
    InMux I__4891 (
            .O(N__22840),
            .I(N__22837));
    LocalMux I__4890 (
            .O(N__22837),
            .I(\Lab_UT.display.dOutP_0_iv_i_2_3 ));
    InMux I__4889 (
            .O(N__22834),
            .I(N__22831));
    LocalMux I__4888 (
            .O(N__22831),
            .I(N__22828));
    Span4Mux_v I__4887 (
            .O(N__22828),
            .I(N__22824));
    InMux I__4886 (
            .O(N__22827),
            .I(N__22821));
    Span4Mux_h I__4885 (
            .O(N__22824),
            .I(N__22815));
    LocalMux I__4884 (
            .O(N__22821),
            .I(N__22815));
    InMux I__4883 (
            .O(N__22820),
            .I(N__22812));
    Odrv4 I__4882 (
            .O(N__22815),
            .I(L3_tx_data_3));
    LocalMux I__4881 (
            .O(N__22812),
            .I(L3_tx_data_3));
    InMux I__4880 (
            .O(N__22807),
            .I(N__22803));
    CascadeMux I__4879 (
            .O(N__22806),
            .I(N__22800));
    LocalMux I__4878 (
            .O(N__22803),
            .I(N__22797));
    InMux I__4877 (
            .O(N__22800),
            .I(N__22794));
    Span4Mux_h I__4876 (
            .O(N__22797),
            .I(N__22787));
    LocalMux I__4875 (
            .O(N__22794),
            .I(N__22787));
    InMux I__4874 (
            .O(N__22793),
            .I(N__22784));
    CascadeMux I__4873 (
            .O(N__22792),
            .I(N__22781));
    Span4Mux_h I__4872 (
            .O(N__22787),
            .I(N__22776));
    LocalMux I__4871 (
            .O(N__22784),
            .I(N__22776));
    InMux I__4870 (
            .O(N__22781),
            .I(N__22773));
    Span4Mux_h I__4869 (
            .O(N__22776),
            .I(N__22770));
    LocalMux I__4868 (
            .O(N__22773),
            .I(\uu2.r_addrZ0Z_5 ));
    Odrv4 I__4867 (
            .O(N__22770),
            .I(\uu2.r_addrZ0Z_5 ));
    InMux I__4866 (
            .O(N__22765),
            .I(N__22761));
    CascadeMux I__4865 (
            .O(N__22764),
            .I(N__22757));
    LocalMux I__4864 (
            .O(N__22761),
            .I(N__22754));
    InMux I__4863 (
            .O(N__22760),
            .I(N__22751));
    InMux I__4862 (
            .O(N__22757),
            .I(N__22748));
    Span4Mux_h I__4861 (
            .O(N__22754),
            .I(N__22745));
    LocalMux I__4860 (
            .O(N__22751),
            .I(\Lab_UT.di_AMones_0 ));
    LocalMux I__4859 (
            .O(N__22748),
            .I(\Lab_UT.di_AMones_0 ));
    Odrv4 I__4858 (
            .O(N__22745),
            .I(\Lab_UT.di_AMones_0 ));
    InMux I__4857 (
            .O(N__22738),
            .I(N__22735));
    LocalMux I__4856 (
            .O(N__22735),
            .I(N__22730));
    InMux I__4855 (
            .O(N__22734),
            .I(N__22727));
    InMux I__4854 (
            .O(N__22733),
            .I(N__22724));
    Span4Mux_v I__4853 (
            .O(N__22730),
            .I(N__22721));
    LocalMux I__4852 (
            .O(N__22727),
            .I(\Lab_UT.di_AMones_2 ));
    LocalMux I__4851 (
            .O(N__22724),
            .I(\Lab_UT.di_AMones_2 ));
    Odrv4 I__4850 (
            .O(N__22721),
            .I(\Lab_UT.di_AMones_2 ));
    InMux I__4849 (
            .O(N__22714),
            .I(N__22702));
    InMux I__4848 (
            .O(N__22713),
            .I(N__22702));
    InMux I__4847 (
            .O(N__22712),
            .I(N__22702));
    InMux I__4846 (
            .O(N__22711),
            .I(N__22702));
    LocalMux I__4845 (
            .O(N__22702),
            .I(N__22699));
    Span4Mux_v I__4844 (
            .O(N__22699),
            .I(N__22696));
    Odrv4 I__4843 (
            .O(N__22696),
            .I(\Lab_UT.ld_enable_AMones ));
    InMux I__4842 (
            .O(N__22693),
            .I(N__22690));
    LocalMux I__4841 (
            .O(N__22690),
            .I(N__22685));
    InMux I__4840 (
            .O(N__22689),
            .I(N__22682));
    InMux I__4839 (
            .O(N__22688),
            .I(N__22679));
    Span4Mux_h I__4838 (
            .O(N__22685),
            .I(N__22676));
    LocalMux I__4837 (
            .O(N__22682),
            .I(\Lab_UT.di_AMones_3 ));
    LocalMux I__4836 (
            .O(N__22679),
            .I(\Lab_UT.di_AMones_3 ));
    Odrv4 I__4835 (
            .O(N__22676),
            .I(\Lab_UT.di_AMones_3 ));
    CascadeMux I__4834 (
            .O(N__22669),
            .I(\Lab_UT.display.N_88_cascade_ ));
    InMux I__4833 (
            .O(N__22666),
            .I(N__22662));
    CascadeMux I__4832 (
            .O(N__22665),
            .I(N__22658));
    LocalMux I__4831 (
            .O(N__22662),
            .I(N__22655));
    InMux I__4830 (
            .O(N__22661),
            .I(N__22652));
    InMux I__4829 (
            .O(N__22658),
            .I(N__22649));
    Odrv12 I__4828 (
            .O(N__22655),
            .I(L3_tx_data_1));
    LocalMux I__4827 (
            .O(N__22652),
            .I(L3_tx_data_1));
    LocalMux I__4826 (
            .O(N__22649),
            .I(L3_tx_data_1));
    CascadeMux I__4825 (
            .O(N__22642),
            .I(\Lab_UT.display.N_120_cascade_ ));
    InMux I__4824 (
            .O(N__22639),
            .I(N__22636));
    LocalMux I__4823 (
            .O(N__22636),
            .I(N__22633));
    Span4Mux_h I__4822 (
            .O(N__22633),
            .I(N__22628));
    InMux I__4821 (
            .O(N__22632),
            .I(N__22623));
    InMux I__4820 (
            .O(N__22631),
            .I(N__22623));
    Odrv4 I__4819 (
            .O(N__22628),
            .I(L3_tx_data_4));
    LocalMux I__4818 (
            .O(N__22623),
            .I(L3_tx_data_4));
    InMux I__4817 (
            .O(N__22618),
            .I(N__22615));
    LocalMux I__4816 (
            .O(N__22615),
            .I(N__22610));
    InMux I__4815 (
            .O(N__22614),
            .I(N__22605));
    InMux I__4814 (
            .O(N__22613),
            .I(N__22605));
    Odrv12 I__4813 (
            .O(N__22610),
            .I(L3_tx_data_5));
    LocalMux I__4812 (
            .O(N__22605),
            .I(L3_tx_data_5));
    CascadeMux I__4811 (
            .O(N__22600),
            .I(\Lab_UT.display.N_153_cascade_ ));
    InMux I__4810 (
            .O(N__22597),
            .I(N__22582));
    InMux I__4809 (
            .O(N__22596),
            .I(N__22582));
    InMux I__4808 (
            .O(N__22595),
            .I(N__22582));
    InMux I__4807 (
            .O(N__22594),
            .I(N__22582));
    InMux I__4806 (
            .O(N__22593),
            .I(N__22582));
    LocalMux I__4805 (
            .O(N__22582),
            .I(\Lab_UT.uu0.l_precountZ0Z_1 ));
    InMux I__4804 (
            .O(N__22579),
            .I(N__22569));
    InMux I__4803 (
            .O(N__22578),
            .I(N__22569));
    InMux I__4802 (
            .O(N__22577),
            .I(N__22569));
    InMux I__4801 (
            .O(N__22576),
            .I(N__22566));
    LocalMux I__4800 (
            .O(N__22569),
            .I(\Lab_UT.uu0.l_countZ0Z_16 ));
    LocalMux I__4799 (
            .O(N__22566),
            .I(\Lab_UT.uu0.l_countZ0Z_16 ));
    CascadeMux I__4798 (
            .O(N__22561),
            .I(N__22557));
    InMux I__4797 (
            .O(N__22560),
            .I(N__22551));
    InMux I__4796 (
            .O(N__22557),
            .I(N__22551));
    InMux I__4795 (
            .O(N__22556),
            .I(N__22548));
    LocalMux I__4794 (
            .O(N__22551),
            .I(N__22543));
    LocalMux I__4793 (
            .O(N__22548),
            .I(N__22543));
    Odrv4 I__4792 (
            .O(N__22543),
            .I(\Lab_UT.uu0.l_countZ0Z_11 ));
    CascadeMux I__4791 (
            .O(N__22540),
            .I(N__22534));
    InMux I__4790 (
            .O(N__22539),
            .I(N__22525));
    InMux I__4789 (
            .O(N__22538),
            .I(N__22525));
    InMux I__4788 (
            .O(N__22537),
            .I(N__22525));
    InMux I__4787 (
            .O(N__22534),
            .I(N__22525));
    LocalMux I__4786 (
            .O(N__22525),
            .I(\Lab_UT.uu0.l_precountZ0Z_2 ));
    CascadeMux I__4785 (
            .O(N__22522),
            .I(N__22516));
    InMux I__4784 (
            .O(N__22521),
            .I(N__22506));
    InMux I__4783 (
            .O(N__22520),
            .I(N__22506));
    InMux I__4782 (
            .O(N__22519),
            .I(N__22506));
    InMux I__4781 (
            .O(N__22516),
            .I(N__22506));
    InMux I__4780 (
            .O(N__22515),
            .I(N__22503));
    LocalMux I__4779 (
            .O(N__22506),
            .I(\Lab_UT.uu0.l_countZ0Z_0 ));
    LocalMux I__4778 (
            .O(N__22503),
            .I(\Lab_UT.uu0.l_countZ0Z_0 ));
    InMux I__4777 (
            .O(N__22498),
            .I(N__22495));
    LocalMux I__4776 (
            .O(N__22495),
            .I(\Lab_UT.uu0.un4_l_count_13 ));
    CascadeMux I__4775 (
            .O(N__22492),
            .I(N__22489));
    InMux I__4774 (
            .O(N__22489),
            .I(N__22481));
    InMux I__4773 (
            .O(N__22488),
            .I(N__22481));
    InMux I__4772 (
            .O(N__22487),
            .I(N__22478));
    InMux I__4771 (
            .O(N__22486),
            .I(N__22475));
    LocalMux I__4770 (
            .O(N__22481),
            .I(N__22472));
    LocalMux I__4769 (
            .O(N__22478),
            .I(N__22469));
    LocalMux I__4768 (
            .O(N__22475),
            .I(\uu2.w_addr_userZ0Z_5 ));
    Odrv12 I__4767 (
            .O(N__22472),
            .I(\uu2.w_addr_userZ0Z_5 ));
    Odrv4 I__4766 (
            .O(N__22469),
            .I(\uu2.w_addr_userZ0Z_5 ));
    CascadeMux I__4765 (
            .O(N__22462),
            .I(N__22456));
    InMux I__4764 (
            .O(N__22461),
            .I(N__22450));
    InMux I__4763 (
            .O(N__22460),
            .I(N__22450));
    InMux I__4762 (
            .O(N__22459),
            .I(N__22447));
    InMux I__4761 (
            .O(N__22456),
            .I(N__22442));
    InMux I__4760 (
            .O(N__22455),
            .I(N__22442));
    LocalMux I__4759 (
            .O(N__22450),
            .I(N__22439));
    LocalMux I__4758 (
            .O(N__22447),
            .I(N__22436));
    LocalMux I__4757 (
            .O(N__22442),
            .I(\uu2.w_addr_userZ0Z_4 ));
    Odrv12 I__4756 (
            .O(N__22439),
            .I(\uu2.w_addr_userZ0Z_4 ));
    Odrv4 I__4755 (
            .O(N__22436),
            .I(\uu2.w_addr_userZ0Z_4 ));
    InMux I__4754 (
            .O(N__22429),
            .I(N__22416));
    InMux I__4753 (
            .O(N__22428),
            .I(N__22416));
    InMux I__4752 (
            .O(N__22427),
            .I(N__22416));
    InMux I__4751 (
            .O(N__22426),
            .I(N__22409));
    InMux I__4750 (
            .O(N__22425),
            .I(N__22409));
    InMux I__4749 (
            .O(N__22424),
            .I(N__22409));
    InMux I__4748 (
            .O(N__22423),
            .I(N__22406));
    LocalMux I__4747 (
            .O(N__22416),
            .I(\uu2.un28_w_addr_user_i ));
    LocalMux I__4746 (
            .O(N__22409),
            .I(\uu2.un28_w_addr_user_i ));
    LocalMux I__4745 (
            .O(N__22406),
            .I(\uu2.un28_w_addr_user_i ));
    InMux I__4744 (
            .O(N__22399),
            .I(N__22390));
    InMux I__4743 (
            .O(N__22398),
            .I(N__22390));
    InMux I__4742 (
            .O(N__22397),
            .I(N__22383));
    InMux I__4741 (
            .O(N__22396),
            .I(N__22383));
    InMux I__4740 (
            .O(N__22395),
            .I(N__22383));
    LocalMux I__4739 (
            .O(N__22390),
            .I(\uu2.un404_ci ));
    LocalMux I__4738 (
            .O(N__22383),
            .I(\uu2.un404_ci ));
    CascadeMux I__4737 (
            .O(N__22378),
            .I(N__22375));
    InMux I__4736 (
            .O(N__22375),
            .I(N__22371));
    CascadeMux I__4735 (
            .O(N__22374),
            .I(N__22367));
    LocalMux I__4734 (
            .O(N__22371),
            .I(N__22364));
    InMux I__4733 (
            .O(N__22370),
            .I(N__22359));
    InMux I__4732 (
            .O(N__22367),
            .I(N__22359));
    Odrv4 I__4731 (
            .O(N__22364),
            .I(\uu2.un426_ci_3 ));
    LocalMux I__4730 (
            .O(N__22359),
            .I(\uu2.un426_ci_3 ));
    InMux I__4729 (
            .O(N__22354),
            .I(N__22343));
    InMux I__4728 (
            .O(N__22353),
            .I(N__22343));
    InMux I__4727 (
            .O(N__22352),
            .I(N__22343));
    InMux I__4726 (
            .O(N__22351),
            .I(N__22340));
    InMux I__4725 (
            .O(N__22350),
            .I(N__22337));
    LocalMux I__4724 (
            .O(N__22343),
            .I(N__22332));
    LocalMux I__4723 (
            .O(N__22340),
            .I(N__22332));
    LocalMux I__4722 (
            .O(N__22337),
            .I(\uu2.w_addr_userZ0Z_6 ));
    Odrv4 I__4721 (
            .O(N__22332),
            .I(\uu2.w_addr_userZ0Z_6 ));
    SRMux I__4720 (
            .O(N__22327),
            .I(N__22323));
    SRMux I__4719 (
            .O(N__22326),
            .I(N__22319));
    LocalMux I__4718 (
            .O(N__22323),
            .I(N__22316));
    SRMux I__4717 (
            .O(N__22322),
            .I(N__22313));
    LocalMux I__4716 (
            .O(N__22319),
            .I(N__22307));
    Span4Mux_h I__4715 (
            .O(N__22316),
            .I(N__22307));
    LocalMux I__4714 (
            .O(N__22313),
            .I(N__22304));
    InMux I__4713 (
            .O(N__22312),
            .I(N__22301));
    Odrv4 I__4712 (
            .O(N__22307),
            .I(\uu2.w_addr_user_RNIMJ3O2Z0Z_2 ));
    Odrv4 I__4711 (
            .O(N__22304),
            .I(\uu2.w_addr_user_RNIMJ3O2Z0Z_2 ));
    LocalMux I__4710 (
            .O(N__22301),
            .I(\uu2.w_addr_user_RNIMJ3O2Z0Z_2 ));
    InMux I__4709 (
            .O(N__22294),
            .I(N__22285));
    InMux I__4708 (
            .O(N__22293),
            .I(N__22285));
    InMux I__4707 (
            .O(N__22292),
            .I(N__22285));
    LocalMux I__4706 (
            .O(N__22285),
            .I(L3_tx_data_rdy));
    CascadeMux I__4705 (
            .O(N__22282),
            .I(N__22277));
    InMux I__4704 (
            .O(N__22281),
            .I(N__22272));
    InMux I__4703 (
            .O(N__22280),
            .I(N__22272));
    InMux I__4702 (
            .O(N__22277),
            .I(N__22269));
    LocalMux I__4701 (
            .O(N__22272),
            .I(L3_tx_data_6));
    LocalMux I__4700 (
            .O(N__22269),
            .I(L3_tx_data_6));
    InMux I__4699 (
            .O(N__22264),
            .I(N__22261));
    LocalMux I__4698 (
            .O(N__22261),
            .I(N__22256));
    InMux I__4697 (
            .O(N__22260),
            .I(N__22251));
    InMux I__4696 (
            .O(N__22259),
            .I(N__22251));
    Span4Mux_h I__4695 (
            .O(N__22256),
            .I(N__22248));
    LocalMux I__4694 (
            .O(N__22251),
            .I(\Lab_UT.uu0.l_countZ0Z_3 ));
    Odrv4 I__4693 (
            .O(N__22248),
            .I(\Lab_UT.uu0.l_countZ0Z_3 ));
    InMux I__4692 (
            .O(N__22243),
            .I(N__22236));
    InMux I__4691 (
            .O(N__22242),
            .I(N__22236));
    InMux I__4690 (
            .O(N__22241),
            .I(N__22232));
    LocalMux I__4689 (
            .O(N__22236),
            .I(N__22229));
    InMux I__4688 (
            .O(N__22235),
            .I(N__22226));
    LocalMux I__4687 (
            .O(N__22232),
            .I(\Lab_UT.uu0.l_countZ0Z_2 ));
    Odrv4 I__4686 (
            .O(N__22229),
            .I(\Lab_UT.uu0.l_countZ0Z_2 ));
    LocalMux I__4685 (
            .O(N__22226),
            .I(\Lab_UT.uu0.l_countZ0Z_2 ));
    CascadeMux I__4684 (
            .O(N__22219),
            .I(\Lab_UT.uu0.un66_ci_cascade_ ));
    InMux I__4683 (
            .O(N__22216),
            .I(N__22208));
    InMux I__4682 (
            .O(N__22215),
            .I(N__22208));
    InMux I__4681 (
            .O(N__22214),
            .I(N__22205));
    InMux I__4680 (
            .O(N__22213),
            .I(N__22202));
    LocalMux I__4679 (
            .O(N__22208),
            .I(\Lab_UT.uu0.l_countZ0Z_4 ));
    LocalMux I__4678 (
            .O(N__22205),
            .I(\Lab_UT.uu0.l_countZ0Z_4 ));
    LocalMux I__4677 (
            .O(N__22202),
            .I(\Lab_UT.uu0.l_countZ0Z_4 ));
    InMux I__4676 (
            .O(N__22195),
            .I(N__22187));
    InMux I__4675 (
            .O(N__22194),
            .I(N__22187));
    InMux I__4674 (
            .O(N__22193),
            .I(N__22184));
    InMux I__4673 (
            .O(N__22192),
            .I(N__22181));
    LocalMux I__4672 (
            .O(N__22187),
            .I(\Lab_UT.uu0.un66_ci ));
    LocalMux I__4671 (
            .O(N__22184),
            .I(\Lab_UT.uu0.un66_ci ));
    LocalMux I__4670 (
            .O(N__22181),
            .I(\Lab_UT.uu0.un66_ci ));
    CEMux I__4669 (
            .O(N__22174),
            .I(N__22159));
    CEMux I__4668 (
            .O(N__22173),
            .I(N__22159));
    CEMux I__4667 (
            .O(N__22172),
            .I(N__22159));
    CEMux I__4666 (
            .O(N__22171),
            .I(N__22159));
    CEMux I__4665 (
            .O(N__22170),
            .I(N__22159));
    GlobalMux I__4664 (
            .O(N__22159),
            .I(N__22156));
    gio2CtrlBuf I__4663 (
            .O(N__22156),
            .I(\Lab_UT.uu0.un11_l_count_i_g ));
    InMux I__4662 (
            .O(N__22153),
            .I(N__22150));
    LocalMux I__4661 (
            .O(N__22150),
            .I(N__22147));
    Span4Mux_v I__4660 (
            .O(N__22147),
            .I(N__22143));
    InMux I__4659 (
            .O(N__22146),
            .I(N__22140));
    Span4Mux_h I__4658 (
            .O(N__22143),
            .I(N__22135));
    LocalMux I__4657 (
            .O(N__22140),
            .I(N__22135));
    Span4Mux_v I__4656 (
            .O(N__22135),
            .I(N__22132));
    Odrv4 I__4655 (
            .O(N__22132),
            .I(\Lab_UT.uu0.delay_lineZ0Z_0 ));
    InMux I__4654 (
            .O(N__22129),
            .I(N__22124));
    InMux I__4653 (
            .O(N__22128),
            .I(N__22121));
    InMux I__4652 (
            .O(N__22127),
            .I(N__22118));
    LocalMux I__4651 (
            .O(N__22124),
            .I(\Lab_UT.uu0.l_countZ0Z_5 ));
    LocalMux I__4650 (
            .O(N__22121),
            .I(\Lab_UT.uu0.l_countZ0Z_5 ));
    LocalMux I__4649 (
            .O(N__22118),
            .I(\Lab_UT.uu0.l_countZ0Z_5 ));
    CascadeMux I__4648 (
            .O(N__22111),
            .I(N__22106));
    CascadeMux I__4647 (
            .O(N__22110),
            .I(N__22103));
    InMux I__4646 (
            .O(N__22109),
            .I(N__22096));
    InMux I__4645 (
            .O(N__22106),
            .I(N__22096));
    InMux I__4644 (
            .O(N__22103),
            .I(N__22096));
    LocalMux I__4643 (
            .O(N__22096),
            .I(\Lab_UT.uu0.l_precountZ0Z_3 ));
    InMux I__4642 (
            .O(N__22093),
            .I(N__22083));
    InMux I__4641 (
            .O(N__22092),
            .I(N__22083));
    InMux I__4640 (
            .O(N__22091),
            .I(N__22083));
    InMux I__4639 (
            .O(N__22090),
            .I(N__22080));
    LocalMux I__4638 (
            .O(N__22083),
            .I(\Lab_UT.uu0.l_countZ0Z_1 ));
    LocalMux I__4637 (
            .O(N__22080),
            .I(\Lab_UT.uu0.l_countZ0Z_1 ));
    InMux I__4636 (
            .O(N__22075),
            .I(N__22072));
    LocalMux I__4635 (
            .O(N__22072),
            .I(N__22068));
    InMux I__4634 (
            .O(N__22071),
            .I(N__22065));
    Span4Mux_h I__4633 (
            .O(N__22068),
            .I(N__22062));
    LocalMux I__4632 (
            .O(N__22065),
            .I(\Lab_UT.uu0.l_countZ0Z_18 ));
    Odrv4 I__4631 (
            .O(N__22062),
            .I(\Lab_UT.uu0.l_countZ0Z_18 ));
    InMux I__4630 (
            .O(N__22057),
            .I(N__22052));
    InMux I__4629 (
            .O(N__22056),
            .I(N__22049));
    InMux I__4628 (
            .O(N__22055),
            .I(N__22046));
    LocalMux I__4627 (
            .O(N__22052),
            .I(\Lab_UT.uu0.l_countZ0Z_15 ));
    LocalMux I__4626 (
            .O(N__22049),
            .I(\Lab_UT.uu0.l_countZ0Z_15 ));
    LocalMux I__4625 (
            .O(N__22046),
            .I(\Lab_UT.uu0.l_countZ0Z_15 ));
    CascadeMux I__4624 (
            .O(N__22039),
            .I(\Lab_UT.uu0.un4_l_count_11_cascade_ ));
    InMux I__4623 (
            .O(N__22036),
            .I(N__22026));
    InMux I__4622 (
            .O(N__22035),
            .I(N__22026));
    InMux I__4621 (
            .O(N__22034),
            .I(N__22026));
    InMux I__4620 (
            .O(N__22033),
            .I(N__22023));
    LocalMux I__4619 (
            .O(N__22026),
            .I(\Lab_UT.uu0.l_countZ0Z_6 ));
    LocalMux I__4618 (
            .O(N__22023),
            .I(\Lab_UT.uu0.l_countZ0Z_6 ));
    InMux I__4617 (
            .O(N__22018),
            .I(N__22015));
    LocalMux I__4616 (
            .O(N__22015),
            .I(N__22012));
    Odrv4 I__4615 (
            .O(N__22012),
            .I(\Lab_UT.uu0.un4_l_count_12 ));
    CascadeMux I__4614 (
            .O(N__22009),
            .I(\Lab_UT.uu0.un4_l_count_16_cascade_ ));
    InMux I__4613 (
            .O(N__22006),
            .I(N__22003));
    LocalMux I__4612 (
            .O(N__22003),
            .I(\Lab_UT.uu0.un4_l_count_18 ));
    InMux I__4611 (
            .O(N__22000),
            .I(N__21996));
    CascadeMux I__4610 (
            .O(N__21999),
            .I(N__21992));
    LocalMux I__4609 (
            .O(N__21996),
            .I(N__21988));
    CascadeMux I__4608 (
            .O(N__21995),
            .I(N__21983));
    InMux I__4607 (
            .O(N__21992),
            .I(N__21980));
    CascadeMux I__4606 (
            .O(N__21991),
            .I(N__21977));
    Span4Mux_v I__4605 (
            .O(N__21988),
            .I(N__21974));
    CascadeMux I__4604 (
            .O(N__21987),
            .I(N__21971));
    InMux I__4603 (
            .O(N__21986),
            .I(N__21966));
    InMux I__4602 (
            .O(N__21983),
            .I(N__21966));
    LocalMux I__4601 (
            .O(N__21980),
            .I(N__21963));
    InMux I__4600 (
            .O(N__21977),
            .I(N__21960));
    Span4Mux_h I__4599 (
            .O(N__21974),
            .I(N__21957));
    InMux I__4598 (
            .O(N__21971),
            .I(N__21954));
    LocalMux I__4597 (
            .O(N__21966),
            .I(N__21949));
    Span4Mux_v I__4596 (
            .O(N__21963),
            .I(N__21949));
    LocalMux I__4595 (
            .O(N__21960),
            .I(N__21946));
    Odrv4 I__4594 (
            .O(N__21957),
            .I(bu_rx_data_6_rep1));
    LocalMux I__4593 (
            .O(N__21954),
            .I(bu_rx_data_6_rep1));
    Odrv4 I__4592 (
            .O(N__21949),
            .I(bu_rx_data_6_rep1));
    Odrv4 I__4591 (
            .O(N__21946),
            .I(bu_rx_data_6_rep1));
    InMux I__4590 (
            .O(N__21937),
            .I(N__21932));
    InMux I__4589 (
            .O(N__21936),
            .I(N__21929));
    InMux I__4588 (
            .O(N__21935),
            .I(N__21926));
    LocalMux I__4587 (
            .O(N__21932),
            .I(N__21919));
    LocalMux I__4586 (
            .O(N__21929),
            .I(N__21919));
    LocalMux I__4585 (
            .O(N__21926),
            .I(N__21915));
    InMux I__4584 (
            .O(N__21925),
            .I(N__21910));
    InMux I__4583 (
            .O(N__21924),
            .I(N__21910));
    Span4Mux_h I__4582 (
            .O(N__21919),
            .I(N__21907));
    InMux I__4581 (
            .O(N__21918),
            .I(N__21904));
    Odrv4 I__4580 (
            .O(N__21915),
            .I(bu_rx_data_5_rep1));
    LocalMux I__4579 (
            .O(N__21910),
            .I(bu_rx_data_5_rep1));
    Odrv4 I__4578 (
            .O(N__21907),
            .I(bu_rx_data_5_rep1));
    LocalMux I__4577 (
            .O(N__21904),
            .I(bu_rx_data_5_rep1));
    InMux I__4576 (
            .O(N__21895),
            .I(N__21892));
    LocalMux I__4575 (
            .O(N__21892),
            .I(N__21888));
    InMux I__4574 (
            .O(N__21891),
            .I(N__21885));
    Span4Mux_h I__4573 (
            .O(N__21888),
            .I(N__21882));
    LocalMux I__4572 (
            .O(N__21885),
            .I(bu_rx_data_fast_3));
    Odrv4 I__4571 (
            .O(N__21882),
            .I(bu_rx_data_fast_3));
    InMux I__4570 (
            .O(N__21877),
            .I(N__21873));
    InMux I__4569 (
            .O(N__21876),
            .I(N__21868));
    LocalMux I__4568 (
            .O(N__21873),
            .I(N__21865));
    InMux I__4567 (
            .O(N__21872),
            .I(N__21862));
    InMux I__4566 (
            .O(N__21871),
            .I(N__21859));
    LocalMux I__4565 (
            .O(N__21868),
            .I(N__21852));
    Span4Mux_v I__4564 (
            .O(N__21865),
            .I(N__21852));
    LocalMux I__4563 (
            .O(N__21862),
            .I(N__21852));
    LocalMux I__4562 (
            .O(N__21859),
            .I(N__21849));
    Span4Mux_h I__4561 (
            .O(N__21852),
            .I(N__21846));
    Odrv12 I__4560 (
            .O(N__21849),
            .I(\buart.Z_rx.hhZ0Z_1 ));
    Odrv4 I__4559 (
            .O(N__21846),
            .I(\buart.Z_rx.hhZ0Z_1 ));
    InMux I__4558 (
            .O(N__21841),
            .I(N__21838));
    LocalMux I__4557 (
            .O(N__21838),
            .I(N__21834));
    InMux I__4556 (
            .O(N__21837),
            .I(N__21828));
    Span4Mux_s3_h I__4555 (
            .O(N__21834),
            .I(N__21825));
    InMux I__4554 (
            .O(N__21833),
            .I(N__21820));
    InMux I__4553 (
            .O(N__21832),
            .I(N__21820));
    CascadeMux I__4552 (
            .O(N__21831),
            .I(N__21816));
    LocalMux I__4551 (
            .O(N__21828),
            .I(N__21813));
    Span4Mux_h I__4550 (
            .O(N__21825),
            .I(N__21810));
    LocalMux I__4549 (
            .O(N__21820),
            .I(N__21807));
    InMux I__4548 (
            .O(N__21819),
            .I(N__21802));
    InMux I__4547 (
            .O(N__21816),
            .I(N__21802));
    Odrv4 I__4546 (
            .O(N__21813),
            .I(bu_rx_data_7_rep1));
    Odrv4 I__4545 (
            .O(N__21810),
            .I(bu_rx_data_7_rep1));
    Odrv4 I__4544 (
            .O(N__21807),
            .I(bu_rx_data_7_rep1));
    LocalMux I__4543 (
            .O(N__21802),
            .I(bu_rx_data_7_rep1));
    InMux I__4542 (
            .O(N__21793),
            .I(N__21790));
    LocalMux I__4541 (
            .O(N__21790),
            .I(N__21787));
    Odrv4 I__4540 (
            .O(N__21787),
            .I(\Lab_UT.uu0.un44_ci ));
    CascadeMux I__4539 (
            .O(N__21784),
            .I(\Lab_UT.uu0.un44_ci_cascade_ ));
    CascadeMux I__4538 (
            .O(N__21781),
            .I(N__21777));
    CascadeMux I__4537 (
            .O(N__21780),
            .I(N__21774));
    InMux I__4536 (
            .O(N__21777),
            .I(N__21771));
    InMux I__4535 (
            .O(N__21774),
            .I(N__21768));
    LocalMux I__4534 (
            .O(N__21771),
            .I(N__21760));
    LocalMux I__4533 (
            .O(N__21768),
            .I(N__21757));
    CascadeMux I__4532 (
            .O(N__21767),
            .I(N__21753));
    CascadeMux I__4531 (
            .O(N__21766),
            .I(N__21750));
    InMux I__4530 (
            .O(N__21765),
            .I(N__21742));
    InMux I__4529 (
            .O(N__21764),
            .I(N__21742));
    InMux I__4528 (
            .O(N__21763),
            .I(N__21742));
    Span4Mux_h I__4527 (
            .O(N__21760),
            .I(N__21739));
    Span4Mux_h I__4526 (
            .O(N__21757),
            .I(N__21736));
    InMux I__4525 (
            .O(N__21756),
            .I(N__21727));
    InMux I__4524 (
            .O(N__21753),
            .I(N__21727));
    InMux I__4523 (
            .O(N__21750),
            .I(N__21727));
    InMux I__4522 (
            .O(N__21749),
            .I(N__21727));
    LocalMux I__4521 (
            .O(N__21742),
            .I(bu_rx_data_3_rep1));
    Odrv4 I__4520 (
            .O(N__21739),
            .I(bu_rx_data_3_rep1));
    Odrv4 I__4519 (
            .O(N__21736),
            .I(bu_rx_data_3_rep1));
    LocalMux I__4518 (
            .O(N__21727),
            .I(bu_rx_data_3_rep1));
    CascadeMux I__4517 (
            .O(N__21718),
            .I(\Lab_UT.dictrl.g1_5_1_cascade_ ));
    InMux I__4516 (
            .O(N__21715),
            .I(N__21712));
    LocalMux I__4515 (
            .O(N__21712),
            .I(N__21709));
    Span4Mux_v I__4514 (
            .O(N__21709),
            .I(N__21706));
    Odrv4 I__4513 (
            .O(N__21706),
            .I(\Lab_UT.dictrl.g1_7_1 ));
    InMux I__4512 (
            .O(N__21703),
            .I(N__21700));
    LocalMux I__4511 (
            .O(N__21700),
            .I(N__21692));
    InMux I__4510 (
            .O(N__21699),
            .I(N__21689));
    CascadeMux I__4509 (
            .O(N__21698),
            .I(N__21686));
    InMux I__4508 (
            .O(N__21697),
            .I(N__21680));
    InMux I__4507 (
            .O(N__21696),
            .I(N__21675));
    InMux I__4506 (
            .O(N__21695),
            .I(N__21675));
    Span4Mux_h I__4505 (
            .O(N__21692),
            .I(N__21672));
    LocalMux I__4504 (
            .O(N__21689),
            .I(N__21669));
    InMux I__4503 (
            .O(N__21686),
            .I(N__21660));
    InMux I__4502 (
            .O(N__21685),
            .I(N__21660));
    InMux I__4501 (
            .O(N__21684),
            .I(N__21660));
    InMux I__4500 (
            .O(N__21683),
            .I(N__21660));
    LocalMux I__4499 (
            .O(N__21680),
            .I(bu_rx_data_2_rep1));
    LocalMux I__4498 (
            .O(N__21675),
            .I(bu_rx_data_2_rep1));
    Odrv4 I__4497 (
            .O(N__21672),
            .I(bu_rx_data_2_rep1));
    Odrv12 I__4496 (
            .O(N__21669),
            .I(bu_rx_data_2_rep1));
    LocalMux I__4495 (
            .O(N__21660),
            .I(bu_rx_data_2_rep1));
    InMux I__4494 (
            .O(N__21649),
            .I(N__21646));
    LocalMux I__4493 (
            .O(N__21646),
            .I(N__21643));
    Odrv4 I__4492 (
            .O(N__21643),
            .I(\Lab_UT.dictrl.g1_4_1 ));
    InMux I__4491 (
            .O(N__21640),
            .I(N__21637));
    LocalMux I__4490 (
            .O(N__21637),
            .I(\Lab_UT.dictrl.currState_fast_3 ));
    InMux I__4489 (
            .O(N__21634),
            .I(N__21631));
    LocalMux I__4488 (
            .O(N__21631),
            .I(N__21628));
    Odrv4 I__4487 (
            .O(N__21628),
            .I(\buart.Z_rx.G_30_0_o3_1_4 ));
    InMux I__4486 (
            .O(N__21625),
            .I(N__21611));
    InMux I__4485 (
            .O(N__21624),
            .I(N__21603));
    InMux I__4484 (
            .O(N__21623),
            .I(N__21598));
    InMux I__4483 (
            .O(N__21622),
            .I(N__21598));
    InMux I__4482 (
            .O(N__21621),
            .I(N__21581));
    InMux I__4481 (
            .O(N__21620),
            .I(N__21581));
    InMux I__4480 (
            .O(N__21619),
            .I(N__21581));
    InMux I__4479 (
            .O(N__21618),
            .I(N__21581));
    InMux I__4478 (
            .O(N__21617),
            .I(N__21581));
    InMux I__4477 (
            .O(N__21616),
            .I(N__21581));
    InMux I__4476 (
            .O(N__21615),
            .I(N__21581));
    InMux I__4475 (
            .O(N__21614),
            .I(N__21581));
    LocalMux I__4474 (
            .O(N__21611),
            .I(N__21578));
    CascadeMux I__4473 (
            .O(N__21610),
            .I(N__21569));
    CascadeMux I__4472 (
            .O(N__21609),
            .I(N__21565));
    InMux I__4471 (
            .O(N__21608),
            .I(N__21562));
    InMux I__4470 (
            .O(N__21607),
            .I(N__21559));
    InMux I__4469 (
            .O(N__21606),
            .I(N__21556));
    LocalMux I__4468 (
            .O(N__21603),
            .I(N__21553));
    LocalMux I__4467 (
            .O(N__21598),
            .I(N__21550));
    LocalMux I__4466 (
            .O(N__21581),
            .I(N__21547));
    Span4Mux_s1_h I__4465 (
            .O(N__21578),
            .I(N__21544));
    InMux I__4464 (
            .O(N__21577),
            .I(N__21537));
    InMux I__4463 (
            .O(N__21576),
            .I(N__21537));
    InMux I__4462 (
            .O(N__21575),
            .I(N__21537));
    InMux I__4461 (
            .O(N__21574),
            .I(N__21529));
    InMux I__4460 (
            .O(N__21573),
            .I(N__21529));
    InMux I__4459 (
            .O(N__21572),
            .I(N__21529));
    InMux I__4458 (
            .O(N__21569),
            .I(N__21522));
    InMux I__4457 (
            .O(N__21568),
            .I(N__21522));
    InMux I__4456 (
            .O(N__21565),
            .I(N__21522));
    LocalMux I__4455 (
            .O(N__21562),
            .I(N__21508));
    LocalMux I__4454 (
            .O(N__21559),
            .I(N__21508));
    LocalMux I__4453 (
            .O(N__21556),
            .I(N__21501));
    Span4Mux_v I__4452 (
            .O(N__21553),
            .I(N__21501));
    Span4Mux_v I__4451 (
            .O(N__21550),
            .I(N__21501));
    Span4Mux_h I__4450 (
            .O(N__21547),
            .I(N__21496));
    Span4Mux_h I__4449 (
            .O(N__21544),
            .I(N__21496));
    LocalMux I__4448 (
            .O(N__21537),
            .I(N__21493));
    InMux I__4447 (
            .O(N__21536),
            .I(N__21490));
    LocalMux I__4446 (
            .O(N__21529),
            .I(N__21485));
    LocalMux I__4445 (
            .O(N__21522),
            .I(N__21485));
    InMux I__4444 (
            .O(N__21521),
            .I(N__21470));
    InMux I__4443 (
            .O(N__21520),
            .I(N__21470));
    InMux I__4442 (
            .O(N__21519),
            .I(N__21470));
    InMux I__4441 (
            .O(N__21518),
            .I(N__21470));
    InMux I__4440 (
            .O(N__21517),
            .I(N__21470));
    InMux I__4439 (
            .O(N__21516),
            .I(N__21470));
    InMux I__4438 (
            .O(N__21515),
            .I(N__21470));
    InMux I__4437 (
            .O(N__21514),
            .I(N__21465));
    InMux I__4436 (
            .O(N__21513),
            .I(N__21465));
    Span4Mux_v I__4435 (
            .O(N__21508),
            .I(N__21462));
    Odrv4 I__4434 (
            .O(N__21501),
            .I(\Lab_UT.dictrl.nextStateZ0Z_3 ));
    Odrv4 I__4433 (
            .O(N__21496),
            .I(\Lab_UT.dictrl.nextStateZ0Z_3 ));
    Odrv12 I__4432 (
            .O(N__21493),
            .I(\Lab_UT.dictrl.nextStateZ0Z_3 ));
    LocalMux I__4431 (
            .O(N__21490),
            .I(\Lab_UT.dictrl.nextStateZ0Z_3 ));
    Odrv4 I__4430 (
            .O(N__21485),
            .I(\Lab_UT.dictrl.nextStateZ0Z_3 ));
    LocalMux I__4429 (
            .O(N__21470),
            .I(\Lab_UT.dictrl.nextStateZ0Z_3 ));
    LocalMux I__4428 (
            .O(N__21465),
            .I(\Lab_UT.dictrl.nextStateZ0Z_3 ));
    Odrv4 I__4427 (
            .O(N__21462),
            .I(\Lab_UT.dictrl.nextStateZ0Z_3 ));
    InMux I__4426 (
            .O(N__21445),
            .I(N__21438));
    InMux I__4425 (
            .O(N__21444),
            .I(N__21435));
    InMux I__4424 (
            .O(N__21443),
            .I(N__21430));
    InMux I__4423 (
            .O(N__21442),
            .I(N__21430));
    InMux I__4422 (
            .O(N__21441),
            .I(N__21427));
    LocalMux I__4421 (
            .O(N__21438),
            .I(N__21420));
    LocalMux I__4420 (
            .O(N__21435),
            .I(N__21420));
    LocalMux I__4419 (
            .O(N__21430),
            .I(N__21420));
    LocalMux I__4418 (
            .O(N__21427),
            .I(bu_rx_data_4_rep1));
    Odrv12 I__4417 (
            .O(N__21420),
            .I(bu_rx_data_4_rep1));
    InMux I__4416 (
            .O(N__21415),
            .I(N__21411));
    InMux I__4415 (
            .O(N__21414),
            .I(N__21408));
    LocalMux I__4414 (
            .O(N__21411),
            .I(N__21403));
    LocalMux I__4413 (
            .O(N__21408),
            .I(N__21400));
    InMux I__4412 (
            .O(N__21407),
            .I(N__21395));
    InMux I__4411 (
            .O(N__21406),
            .I(N__21395));
    Span4Mux_v I__4410 (
            .O(N__21403),
            .I(N__21384));
    Span4Mux_s2_v I__4409 (
            .O(N__21400),
            .I(N__21384));
    LocalMux I__4408 (
            .O(N__21395),
            .I(N__21381));
    InMux I__4407 (
            .O(N__21394),
            .I(N__21376));
    InMux I__4406 (
            .O(N__21393),
            .I(N__21376));
    InMux I__4405 (
            .O(N__21392),
            .I(N__21367));
    InMux I__4404 (
            .O(N__21391),
            .I(N__21367));
    InMux I__4403 (
            .O(N__21390),
            .I(N__21367));
    InMux I__4402 (
            .O(N__21389),
            .I(N__21367));
    Odrv4 I__4401 (
            .O(N__21384),
            .I(bu_rx_data_1_rep1));
    Odrv12 I__4400 (
            .O(N__21381),
            .I(bu_rx_data_1_rep1));
    LocalMux I__4399 (
            .O(N__21376),
            .I(bu_rx_data_1_rep1));
    LocalMux I__4398 (
            .O(N__21367),
            .I(bu_rx_data_1_rep1));
    InMux I__4397 (
            .O(N__21358),
            .I(N__21355));
    LocalMux I__4396 (
            .O(N__21355),
            .I(\Lab_UT.dictrl.decoder.g0Z0Z_3 ));
    InMux I__4395 (
            .O(N__21352),
            .I(N__21348));
    InMux I__4394 (
            .O(N__21351),
            .I(N__21343));
    LocalMux I__4393 (
            .O(N__21348),
            .I(N__21340));
    InMux I__4392 (
            .O(N__21347),
            .I(N__21335));
    InMux I__4391 (
            .O(N__21346),
            .I(N__21335));
    LocalMux I__4390 (
            .O(N__21343),
            .I(N__21330));
    Span4Mux_v I__4389 (
            .O(N__21340),
            .I(N__21330));
    LocalMux I__4388 (
            .O(N__21335),
            .I(bu_rx_data_0_rep1));
    Odrv4 I__4387 (
            .O(N__21330),
            .I(bu_rx_data_0_rep1));
    InMux I__4386 (
            .O(N__21325),
            .I(N__21322));
    LocalMux I__4385 (
            .O(N__21322),
            .I(\Lab_UT.dictrl.r_dicLdMtens14_i_6 ));
    InMux I__4384 (
            .O(N__21319),
            .I(N__21316));
    LocalMux I__4383 (
            .O(N__21316),
            .I(N__21313));
    Span4Mux_h I__4382 (
            .O(N__21313),
            .I(N__21310));
    Odrv4 I__4381 (
            .O(N__21310),
            .I(\Lab_UT.dictrl.r_dicLdMtens20_i_6 ));
    InMux I__4380 (
            .O(N__21307),
            .I(N__21304));
    LocalMux I__4379 (
            .O(N__21304),
            .I(N__21301));
    Span4Mux_h I__4378 (
            .O(N__21301),
            .I(N__21298));
    Odrv4 I__4377 (
            .O(N__21298),
            .I(\Lab_UT.dictrl.r_enable3_3_iv_1 ));
    CascadeMux I__4376 (
            .O(N__21295),
            .I(\buart.Z_rx.G_30_0_o3_1_0_cascade_ ));
    InMux I__4375 (
            .O(N__21292),
            .I(N__21287));
    InMux I__4374 (
            .O(N__21291),
            .I(N__21281));
    InMux I__4373 (
            .O(N__21290),
            .I(N__21281));
    LocalMux I__4372 (
            .O(N__21287),
            .I(N__21278));
    InMux I__4371 (
            .O(N__21286),
            .I(N__21275));
    LocalMux I__4370 (
            .O(N__21281),
            .I(Lab_UT_dictrl_decoder_de_cr_1));
    Odrv4 I__4369 (
            .O(N__21278),
            .I(Lab_UT_dictrl_decoder_de_cr_1));
    LocalMux I__4368 (
            .O(N__21275),
            .I(Lab_UT_dictrl_decoder_de_cr_1));
    CascadeMux I__4367 (
            .O(N__21268),
            .I(N__21261));
    InMux I__4366 (
            .O(N__21267),
            .I(N__21254));
    InMux I__4365 (
            .O(N__21266),
            .I(N__21254));
    CascadeMux I__4364 (
            .O(N__21265),
            .I(N__21251));
    CascadeMux I__4363 (
            .O(N__21264),
            .I(N__21247));
    InMux I__4362 (
            .O(N__21261),
            .I(N__21241));
    InMux I__4361 (
            .O(N__21260),
            .I(N__21238));
    InMux I__4360 (
            .O(N__21259),
            .I(N__21235));
    LocalMux I__4359 (
            .O(N__21254),
            .I(N__21231));
    InMux I__4358 (
            .O(N__21251),
            .I(N__21228));
    InMux I__4357 (
            .O(N__21250),
            .I(N__21223));
    InMux I__4356 (
            .O(N__21247),
            .I(N__21223));
    InMux I__4355 (
            .O(N__21246),
            .I(N__21219));
    InMux I__4354 (
            .O(N__21245),
            .I(N__21215));
    CascadeMux I__4353 (
            .O(N__21244),
            .I(N__21212));
    LocalMux I__4352 (
            .O(N__21241),
            .I(N__21207));
    LocalMux I__4351 (
            .O(N__21238),
            .I(N__21207));
    LocalMux I__4350 (
            .O(N__21235),
            .I(N__21204));
    InMux I__4349 (
            .O(N__21234),
            .I(N__21201));
    Span4Mux_v I__4348 (
            .O(N__21231),
            .I(N__21194));
    LocalMux I__4347 (
            .O(N__21228),
            .I(N__21194));
    LocalMux I__4346 (
            .O(N__21223),
            .I(N__21194));
    InMux I__4345 (
            .O(N__21222),
            .I(N__21191));
    LocalMux I__4344 (
            .O(N__21219),
            .I(N__21188));
    InMux I__4343 (
            .O(N__21218),
            .I(N__21185));
    LocalMux I__4342 (
            .O(N__21215),
            .I(N__21182));
    InMux I__4341 (
            .O(N__21212),
            .I(N__21179));
    Span4Mux_v I__4340 (
            .O(N__21207),
            .I(N__21176));
    Span4Mux_h I__4339 (
            .O(N__21204),
            .I(N__21171));
    LocalMux I__4338 (
            .O(N__21201),
            .I(N__21171));
    Span4Mux_v I__4337 (
            .O(N__21194),
            .I(N__21168));
    LocalMux I__4336 (
            .O(N__21191),
            .I(N__21165));
    Span4Mux_v I__4335 (
            .O(N__21188),
            .I(N__21160));
    LocalMux I__4334 (
            .O(N__21185),
            .I(N__21160));
    Span4Mux_s3_h I__4333 (
            .O(N__21182),
            .I(N__21157));
    LocalMux I__4332 (
            .O(N__21179),
            .I(N__21152));
    Span4Mux_h I__4331 (
            .O(N__21176),
            .I(N__21152));
    Span4Mux_v I__4330 (
            .O(N__21171),
            .I(N__21147));
    Span4Mux_h I__4329 (
            .O(N__21168),
            .I(N__21147));
    Odrv12 I__4328 (
            .O(N__21165),
            .I(\Lab_UT.dictrl.currStateZ0Z_0 ));
    Odrv4 I__4327 (
            .O(N__21160),
            .I(\Lab_UT.dictrl.currStateZ0Z_0 ));
    Odrv4 I__4326 (
            .O(N__21157),
            .I(\Lab_UT.dictrl.currStateZ0Z_0 ));
    Odrv4 I__4325 (
            .O(N__21152),
            .I(\Lab_UT.dictrl.currStateZ0Z_0 ));
    Odrv4 I__4324 (
            .O(N__21147),
            .I(\Lab_UT.dictrl.currStateZ0Z_0 ));
    CascadeMux I__4323 (
            .O(N__21136),
            .I(N_6_cascade_));
    InMux I__4322 (
            .O(N__21133),
            .I(N__21130));
    LocalMux I__4321 (
            .O(N__21130),
            .I(N__21127));
    Span4Mux_s3_h I__4320 (
            .O(N__21127),
            .I(N__21124));
    Span4Mux_h I__4319 (
            .O(N__21124),
            .I(N__21121));
    Odrv4 I__4318 (
            .O(N__21121),
            .I(\Lab_UT.dictrl.N_21_0 ));
    InMux I__4317 (
            .O(N__21118),
            .I(N__21115));
    LocalMux I__4316 (
            .O(N__21115),
            .I(\resetGen.escKey_4_0 ));
    InMux I__4315 (
            .O(N__21112),
            .I(N__21104));
    InMux I__4314 (
            .O(N__21111),
            .I(N__21099));
    InMux I__4313 (
            .O(N__21110),
            .I(N__21099));
    InMux I__4312 (
            .O(N__21109),
            .I(N__21087));
    InMux I__4311 (
            .O(N__21108),
            .I(N__21084));
    InMux I__4310 (
            .O(N__21107),
            .I(N__21081));
    LocalMux I__4309 (
            .O(N__21104),
            .I(N__21076));
    LocalMux I__4308 (
            .O(N__21099),
            .I(N__21076));
    InMux I__4307 (
            .O(N__21098),
            .I(N__21073));
    InMux I__4306 (
            .O(N__21097),
            .I(N__21054));
    InMux I__4305 (
            .O(N__21096),
            .I(N__21054));
    InMux I__4304 (
            .O(N__21095),
            .I(N__21054));
    InMux I__4303 (
            .O(N__21094),
            .I(N__21054));
    InMux I__4302 (
            .O(N__21093),
            .I(N__21054));
    InMux I__4301 (
            .O(N__21092),
            .I(N__21054));
    InMux I__4300 (
            .O(N__21091),
            .I(N__21054));
    InMux I__4299 (
            .O(N__21090),
            .I(N__21054));
    LocalMux I__4298 (
            .O(N__21087),
            .I(N__21051));
    LocalMux I__4297 (
            .O(N__21084),
            .I(N__21048));
    LocalMux I__4296 (
            .O(N__21081),
            .I(N__21045));
    Span4Mux_v I__4295 (
            .O(N__21076),
            .I(N__21023));
    LocalMux I__4294 (
            .O(N__21073),
            .I(N__21023));
    InMux I__4293 (
            .O(N__21072),
            .I(N__21020));
    InMux I__4292 (
            .O(N__21071),
            .I(N__21017));
    LocalMux I__4291 (
            .O(N__21054),
            .I(N__21008));
    Span4Mux_h I__4290 (
            .O(N__21051),
            .I(N__21008));
    Span4Mux_v I__4289 (
            .O(N__21048),
            .I(N__21008));
    Span4Mux_v I__4288 (
            .O(N__21045),
            .I(N__21008));
    InMux I__4287 (
            .O(N__21044),
            .I(N__21001));
    InMux I__4286 (
            .O(N__21043),
            .I(N__21001));
    InMux I__4285 (
            .O(N__21042),
            .I(N__21001));
    InMux I__4284 (
            .O(N__21041),
            .I(N__20990));
    InMux I__4283 (
            .O(N__21040),
            .I(N__20990));
    InMux I__4282 (
            .O(N__21039),
            .I(N__20990));
    InMux I__4281 (
            .O(N__21038),
            .I(N__20990));
    InMux I__4280 (
            .O(N__21037),
            .I(N__20990));
    InMux I__4279 (
            .O(N__21036),
            .I(N__20985));
    InMux I__4278 (
            .O(N__21035),
            .I(N__20985));
    InMux I__4277 (
            .O(N__21034),
            .I(N__20970));
    InMux I__4276 (
            .O(N__21033),
            .I(N__20970));
    InMux I__4275 (
            .O(N__21032),
            .I(N__20970));
    InMux I__4274 (
            .O(N__21031),
            .I(N__20970));
    InMux I__4273 (
            .O(N__21030),
            .I(N__20970));
    InMux I__4272 (
            .O(N__21029),
            .I(N__20970));
    InMux I__4271 (
            .O(N__21028),
            .I(N__20970));
    Span4Mux_h I__4270 (
            .O(N__21023),
            .I(N__20967));
    LocalMux I__4269 (
            .O(N__21020),
            .I(\Lab_UT.dictrl.nextStateZ0Z_0 ));
    LocalMux I__4268 (
            .O(N__21017),
            .I(\Lab_UT.dictrl.nextStateZ0Z_0 ));
    Odrv4 I__4267 (
            .O(N__21008),
            .I(\Lab_UT.dictrl.nextStateZ0Z_0 ));
    LocalMux I__4266 (
            .O(N__21001),
            .I(\Lab_UT.dictrl.nextStateZ0Z_0 ));
    LocalMux I__4265 (
            .O(N__20990),
            .I(\Lab_UT.dictrl.nextStateZ0Z_0 ));
    LocalMux I__4264 (
            .O(N__20985),
            .I(\Lab_UT.dictrl.nextStateZ0Z_0 ));
    LocalMux I__4263 (
            .O(N__20970),
            .I(\Lab_UT.dictrl.nextStateZ0Z_0 ));
    Odrv4 I__4262 (
            .O(N__20967),
            .I(\Lab_UT.dictrl.nextStateZ0Z_0 ));
    CascadeMux I__4261 (
            .O(N__20950),
            .I(N__20946));
    InMux I__4260 (
            .O(N__20949),
            .I(N__20941));
    InMux I__4259 (
            .O(N__20946),
            .I(N__20941));
    LocalMux I__4258 (
            .O(N__20941),
            .I(N__20932));
    CascadeMux I__4257 (
            .O(N__20940),
            .I(N__20929));
    CascadeMux I__4256 (
            .O(N__20939),
            .I(N__20926));
    InMux I__4255 (
            .O(N__20938),
            .I(N__20923));
    InMux I__4254 (
            .O(N__20937),
            .I(N__20916));
    InMux I__4253 (
            .O(N__20936),
            .I(N__20916));
    InMux I__4252 (
            .O(N__20935),
            .I(N__20916));
    Span4Mux_h I__4251 (
            .O(N__20932),
            .I(N__20913));
    InMux I__4250 (
            .O(N__20929),
            .I(N__20910));
    InMux I__4249 (
            .O(N__20926),
            .I(N__20907));
    LocalMux I__4248 (
            .O(N__20923),
            .I(N__20904));
    LocalMux I__4247 (
            .O(N__20916),
            .I(N__20901));
    Span4Mux_v I__4246 (
            .O(N__20913),
            .I(N__20895));
    LocalMux I__4245 (
            .O(N__20910),
            .I(N__20895));
    LocalMux I__4244 (
            .O(N__20907),
            .I(N__20892));
    Span4Mux_v I__4243 (
            .O(N__20904),
            .I(N__20886));
    Span4Mux_h I__4242 (
            .O(N__20901),
            .I(N__20886));
    InMux I__4241 (
            .O(N__20900),
            .I(N__20883));
    Span4Mux_h I__4240 (
            .O(N__20895),
            .I(N__20880));
    Span4Mux_h I__4239 (
            .O(N__20892),
            .I(N__20877));
    InMux I__4238 (
            .O(N__20891),
            .I(N__20874));
    Span4Mux_h I__4237 (
            .O(N__20886),
            .I(N__20871));
    LocalMux I__4236 (
            .O(N__20883),
            .I(\Lab_UT.dictrl.currState_0_rep2 ));
    Odrv4 I__4235 (
            .O(N__20880),
            .I(\Lab_UT.dictrl.currState_0_rep2 ));
    Odrv4 I__4234 (
            .O(N__20877),
            .I(\Lab_UT.dictrl.currState_0_rep2 ));
    LocalMux I__4233 (
            .O(N__20874),
            .I(\Lab_UT.dictrl.currState_0_rep2 ));
    Odrv4 I__4232 (
            .O(N__20871),
            .I(\Lab_UT.dictrl.currState_0_rep2 ));
    CascadeMux I__4231 (
            .O(N__20860),
            .I(\Lab_UT.dictrl.g0_7_cascade_ ));
    CascadeMux I__4230 (
            .O(N__20857),
            .I(N__20854));
    InMux I__4229 (
            .O(N__20854),
            .I(N__20851));
    LocalMux I__4228 (
            .O(N__20851),
            .I(N__20848));
    Span4Mux_h I__4227 (
            .O(N__20848),
            .I(N__20845));
    Span4Mux_v I__4226 (
            .O(N__20845),
            .I(N__20842));
    Odrv4 I__4225 (
            .O(N__20842),
            .I(\Lab_UT.dictrl.g0_10 ));
    InMux I__4224 (
            .O(N__20839),
            .I(N__20835));
    InMux I__4223 (
            .O(N__20838),
            .I(N__20832));
    LocalMux I__4222 (
            .O(N__20835),
            .I(N__20829));
    LocalMux I__4221 (
            .O(N__20832),
            .I(bu_rx_data_fast_1));
    Odrv4 I__4220 (
            .O(N__20829),
            .I(bu_rx_data_fast_1));
    InMux I__4219 (
            .O(N__20824),
            .I(N__20821));
    LocalMux I__4218 (
            .O(N__20821),
            .I(N__20818));
    Odrv12 I__4217 (
            .O(N__20818),
            .I(\Lab_UT.dictrl.r_dicLdMtens16 ));
    CascadeMux I__4216 (
            .O(N__20815),
            .I(N__20802));
    InMux I__4215 (
            .O(N__20814),
            .I(N__20799));
    InMux I__4214 (
            .O(N__20813),
            .I(N__20796));
    CascadeMux I__4213 (
            .O(N__20812),
            .I(N__20789));
    CascadeMux I__4212 (
            .O(N__20811),
            .I(N__20786));
    CascadeMux I__4211 (
            .O(N__20810),
            .I(N__20783));
    CascadeMux I__4210 (
            .O(N__20809),
            .I(N__20780));
    CascadeMux I__4209 (
            .O(N__20808),
            .I(N__20777));
    CascadeMux I__4208 (
            .O(N__20807),
            .I(N__20774));
    CascadeMux I__4207 (
            .O(N__20806),
            .I(N__20771));
    CascadeMux I__4206 (
            .O(N__20805),
            .I(N__20768));
    InMux I__4205 (
            .O(N__20802),
            .I(N__20764));
    LocalMux I__4204 (
            .O(N__20799),
            .I(N__20761));
    LocalMux I__4203 (
            .O(N__20796),
            .I(N__20758));
    CascadeMux I__4202 (
            .O(N__20795),
            .I(N__20752));
    CascadeMux I__4201 (
            .O(N__20794),
            .I(N__20748));
    CascadeMux I__4200 (
            .O(N__20793),
            .I(N__20743));
    CascadeMux I__4199 (
            .O(N__20792),
            .I(N__20739));
    InMux I__4198 (
            .O(N__20789),
            .I(N__20730));
    InMux I__4197 (
            .O(N__20786),
            .I(N__20730));
    InMux I__4196 (
            .O(N__20783),
            .I(N__20730));
    InMux I__4195 (
            .O(N__20780),
            .I(N__20730));
    InMux I__4194 (
            .O(N__20777),
            .I(N__20721));
    InMux I__4193 (
            .O(N__20774),
            .I(N__20721));
    InMux I__4192 (
            .O(N__20771),
            .I(N__20721));
    InMux I__4191 (
            .O(N__20768),
            .I(N__20721));
    InMux I__4190 (
            .O(N__20767),
            .I(N__20718));
    LocalMux I__4189 (
            .O(N__20764),
            .I(N__20713));
    Span4Mux_h I__4188 (
            .O(N__20761),
            .I(N__20713));
    Span12Mux_s6_h I__4187 (
            .O(N__20758),
            .I(N__20710));
    InMux I__4186 (
            .O(N__20757),
            .I(N__20705));
    InMux I__4185 (
            .O(N__20756),
            .I(N__20705));
    InMux I__4184 (
            .O(N__20755),
            .I(N__20698));
    InMux I__4183 (
            .O(N__20752),
            .I(N__20698));
    InMux I__4182 (
            .O(N__20751),
            .I(N__20698));
    InMux I__4181 (
            .O(N__20748),
            .I(N__20685));
    InMux I__4180 (
            .O(N__20747),
            .I(N__20685));
    InMux I__4179 (
            .O(N__20746),
            .I(N__20685));
    InMux I__4178 (
            .O(N__20743),
            .I(N__20685));
    InMux I__4177 (
            .O(N__20742),
            .I(N__20685));
    InMux I__4176 (
            .O(N__20739),
            .I(N__20685));
    LocalMux I__4175 (
            .O(N__20730),
            .I(\Lab_UT.dictrl.nextStateZ0Z_2 ));
    LocalMux I__4174 (
            .O(N__20721),
            .I(\Lab_UT.dictrl.nextStateZ0Z_2 ));
    LocalMux I__4173 (
            .O(N__20718),
            .I(\Lab_UT.dictrl.nextStateZ0Z_2 ));
    Odrv4 I__4172 (
            .O(N__20713),
            .I(\Lab_UT.dictrl.nextStateZ0Z_2 ));
    Odrv12 I__4171 (
            .O(N__20710),
            .I(\Lab_UT.dictrl.nextStateZ0Z_2 ));
    LocalMux I__4170 (
            .O(N__20705),
            .I(\Lab_UT.dictrl.nextStateZ0Z_2 ));
    LocalMux I__4169 (
            .O(N__20698),
            .I(\Lab_UT.dictrl.nextStateZ0Z_2 ));
    LocalMux I__4168 (
            .O(N__20685),
            .I(\Lab_UT.dictrl.nextStateZ0Z_2 ));
    InMux I__4167 (
            .O(N__20668),
            .I(N__20654));
    InMux I__4166 (
            .O(N__20667),
            .I(N__20644));
    InMux I__4165 (
            .O(N__20666),
            .I(N__20644));
    InMux I__4164 (
            .O(N__20665),
            .I(N__20644));
    InMux I__4163 (
            .O(N__20664),
            .I(N__20644));
    InMux I__4162 (
            .O(N__20663),
            .I(N__20635));
    InMux I__4161 (
            .O(N__20662),
            .I(N__20635));
    InMux I__4160 (
            .O(N__20661),
            .I(N__20635));
    InMux I__4159 (
            .O(N__20660),
            .I(N__20635));
    CascadeMux I__4158 (
            .O(N__20659),
            .I(N__20631));
    CascadeMux I__4157 (
            .O(N__20658),
            .I(N__20628));
    CascadeMux I__4156 (
            .O(N__20657),
            .I(N__20624));
    LocalMux I__4155 (
            .O(N__20654),
            .I(N__20619));
    InMux I__4154 (
            .O(N__20653),
            .I(N__20616));
    LocalMux I__4153 (
            .O(N__20644),
            .I(N__20611));
    LocalMux I__4152 (
            .O(N__20635),
            .I(N__20611));
    InMux I__4151 (
            .O(N__20634),
            .I(N__20598));
    InMux I__4150 (
            .O(N__20631),
            .I(N__20598));
    InMux I__4149 (
            .O(N__20628),
            .I(N__20598));
    InMux I__4148 (
            .O(N__20627),
            .I(N__20598));
    InMux I__4147 (
            .O(N__20624),
            .I(N__20598));
    InMux I__4146 (
            .O(N__20623),
            .I(N__20598));
    InMux I__4145 (
            .O(N__20622),
            .I(N__20595));
    Span4Mux_h I__4144 (
            .O(N__20619),
            .I(N__20592));
    LocalMux I__4143 (
            .O(N__20616),
            .I(N__20585));
    Span12Mux_s6_v I__4142 (
            .O(N__20611),
            .I(N__20585));
    LocalMux I__4141 (
            .O(N__20598),
            .I(N__20585));
    LocalMux I__4140 (
            .O(N__20595),
            .I(\Lab_UT.dictrl.nextStateZ0Z_1 ));
    Odrv4 I__4139 (
            .O(N__20592),
            .I(\Lab_UT.dictrl.nextStateZ0Z_1 ));
    Odrv12 I__4138 (
            .O(N__20585),
            .I(\Lab_UT.dictrl.nextStateZ0Z_1 ));
    InMux I__4137 (
            .O(N__20578),
            .I(N__20575));
    LocalMux I__4136 (
            .O(N__20575),
            .I(N__20572));
    Odrv4 I__4135 (
            .O(N__20572),
            .I(\Lab_UT.dictrl.r_dicLdMtens17 ));
    InMux I__4134 (
            .O(N__20569),
            .I(N__20566));
    LocalMux I__4133 (
            .O(N__20566),
            .I(N__20563));
    Span4Mux_h I__4132 (
            .O(N__20563),
            .I(N__20557));
    InMux I__4131 (
            .O(N__20562),
            .I(N__20554));
    InMux I__4130 (
            .O(N__20561),
            .I(N__20551));
    InMux I__4129 (
            .O(N__20560),
            .I(N__20548));
    Odrv4 I__4128 (
            .O(N__20557),
            .I(\Lab_UT.dictrl.currState_ret_1and ));
    LocalMux I__4127 (
            .O(N__20554),
            .I(\Lab_UT.dictrl.currState_ret_1and ));
    LocalMux I__4126 (
            .O(N__20551),
            .I(\Lab_UT.dictrl.currState_ret_1and ));
    LocalMux I__4125 (
            .O(N__20548),
            .I(\Lab_UT.dictrl.currState_ret_1and ));
    CascadeMux I__4124 (
            .O(N__20539),
            .I(N__20536));
    InMux I__4123 (
            .O(N__20536),
            .I(N__20533));
    LocalMux I__4122 (
            .O(N__20533),
            .I(\Lab_UT.dictrl.dicLdAMones_rst ));
    InMux I__4121 (
            .O(N__20530),
            .I(N__20524));
    InMux I__4120 (
            .O(N__20529),
            .I(N__20524));
    LocalMux I__4119 (
            .O(N__20524),
            .I(\Lab_UT.dictrl.dicLdAMonesZ0 ));
    CascadeMux I__4118 (
            .O(N__20521),
            .I(\Lab_UT.dictrl.dicLdAMones_rst_cascade_ ));
    InMux I__4117 (
            .O(N__20518),
            .I(N__20508));
    InMux I__4116 (
            .O(N__20517),
            .I(N__20508));
    InMux I__4115 (
            .O(N__20516),
            .I(N__20508));
    InMux I__4114 (
            .O(N__20515),
            .I(N__20503));
    LocalMux I__4113 (
            .O(N__20508),
            .I(N__20500));
    InMux I__4112 (
            .O(N__20507),
            .I(N__20495));
    InMux I__4111 (
            .O(N__20506),
            .I(N__20495));
    LocalMux I__4110 (
            .O(N__20503),
            .I(N__20492));
    Span4Mux_h I__4109 (
            .O(N__20500),
            .I(N__20487));
    LocalMux I__4108 (
            .O(N__20495),
            .I(N__20487));
    Span4Mux_v I__4107 (
            .O(N__20492),
            .I(N__20484));
    Span4Mux_v I__4106 (
            .O(N__20487),
            .I(N__20481));
    Odrv4 I__4105 (
            .O(N__20484),
            .I(\Lab_UT.dictrl.r_dicLdMtens23_2 ));
    Odrv4 I__4104 (
            .O(N__20481),
            .I(\Lab_UT.dictrl.r_dicLdMtens23_2 ));
    CascadeMux I__4103 (
            .O(N__20476),
            .I(N__20472));
    InMux I__4102 (
            .O(N__20475),
            .I(N__20469));
    InMux I__4101 (
            .O(N__20472),
            .I(N__20466));
    LocalMux I__4100 (
            .O(N__20469),
            .I(N__20463));
    LocalMux I__4099 (
            .O(N__20466),
            .I(\Lab_UT.dictrl.dicLdAStensZ0 ));
    Odrv12 I__4098 (
            .O(N__20463),
            .I(\Lab_UT.dictrl.dicLdAStensZ0 ));
    InMux I__4097 (
            .O(N__20458),
            .I(N__20454));
    InMux I__4096 (
            .O(N__20457),
            .I(N__20451));
    LocalMux I__4095 (
            .O(N__20454),
            .I(N__20448));
    LocalMux I__4094 (
            .O(N__20451),
            .I(N__20445));
    Span4Mux_v I__4093 (
            .O(N__20448),
            .I(N__20442));
    Span4Mux_v I__4092 (
            .O(N__20445),
            .I(N__20437));
    Span4Mux_h I__4091 (
            .O(N__20442),
            .I(N__20437));
    Odrv4 I__4090 (
            .O(N__20437),
            .I(\Lab_UT.dictrl.dicLdAStens_rst ));
    InMux I__4089 (
            .O(N__20434),
            .I(N__20428));
    InMux I__4088 (
            .O(N__20433),
            .I(N__20428));
    LocalMux I__4087 (
            .O(N__20428),
            .I(N__20425));
    Span4Mux_v I__4086 (
            .O(N__20425),
            .I(N__20419));
    InMux I__4085 (
            .O(N__20424),
            .I(N__20412));
    InMux I__4084 (
            .O(N__20423),
            .I(N__20412));
    InMux I__4083 (
            .O(N__20422),
            .I(N__20412));
    Sp12to4 I__4082 (
            .O(N__20419),
            .I(N__20409));
    LocalMux I__4081 (
            .O(N__20412),
            .I(N__20406));
    Span12Mux_s7_h I__4080 (
            .O(N__20409),
            .I(N__20401));
    Span12Mux_s4_v I__4079 (
            .O(N__20406),
            .I(N__20401));
    Odrv12 I__4078 (
            .O(N__20401),
            .I(\resetGen.escKeyZ0 ));
    CascadeMux I__4077 (
            .O(N__20398),
            .I(N__20389));
    CascadeMux I__4076 (
            .O(N__20397),
            .I(N__20385));
    CascadeMux I__4075 (
            .O(N__20396),
            .I(N__20382));
    InMux I__4074 (
            .O(N__20395),
            .I(N__20379));
    InMux I__4073 (
            .O(N__20394),
            .I(N__20374));
    InMux I__4072 (
            .O(N__20393),
            .I(N__20374));
    InMux I__4071 (
            .O(N__20392),
            .I(N__20371));
    InMux I__4070 (
            .O(N__20389),
            .I(N__20362));
    InMux I__4069 (
            .O(N__20388),
            .I(N__20362));
    InMux I__4068 (
            .O(N__20385),
            .I(N__20362));
    InMux I__4067 (
            .O(N__20382),
            .I(N__20357));
    LocalMux I__4066 (
            .O(N__20379),
            .I(N__20352));
    LocalMux I__4065 (
            .O(N__20374),
            .I(N__20352));
    LocalMux I__4064 (
            .O(N__20371),
            .I(N__20349));
    InMux I__4063 (
            .O(N__20370),
            .I(N__20346));
    InMux I__4062 (
            .O(N__20369),
            .I(N__20343));
    LocalMux I__4061 (
            .O(N__20362),
            .I(N__20340));
    InMux I__4060 (
            .O(N__20361),
            .I(N__20335));
    InMux I__4059 (
            .O(N__20360),
            .I(N__20335));
    LocalMux I__4058 (
            .O(N__20357),
            .I(N__20329));
    Span4Mux_v I__4057 (
            .O(N__20352),
            .I(N__20329));
    Span4Mux_v I__4056 (
            .O(N__20349),
            .I(N__20324));
    LocalMux I__4055 (
            .O(N__20346),
            .I(N__20324));
    LocalMux I__4054 (
            .O(N__20343),
            .I(N__20321));
    Span4Mux_h I__4053 (
            .O(N__20340),
            .I(N__20316));
    LocalMux I__4052 (
            .O(N__20335),
            .I(N__20316));
    InMux I__4051 (
            .O(N__20334),
            .I(N__20313));
    Span4Mux_h I__4050 (
            .O(N__20329),
            .I(N__20308));
    Span4Mux_v I__4049 (
            .O(N__20324),
            .I(N__20308));
    Odrv4 I__4048 (
            .O(N__20321),
            .I(\Lab_UT.dictrl.currState_3_rep1 ));
    Odrv4 I__4047 (
            .O(N__20316),
            .I(\Lab_UT.dictrl.currState_3_rep1 ));
    LocalMux I__4046 (
            .O(N__20313),
            .I(\Lab_UT.dictrl.currState_3_rep1 ));
    Odrv4 I__4045 (
            .O(N__20308),
            .I(\Lab_UT.dictrl.currState_3_rep1 ));
    InMux I__4044 (
            .O(N__20299),
            .I(N__20296));
    LocalMux I__4043 (
            .O(N__20296),
            .I(N__20292));
    InMux I__4042 (
            .O(N__20295),
            .I(N__20289));
    Odrv12 I__4041 (
            .O(N__20292),
            .I(\Lab_UT.dictrl.N_5 ));
    LocalMux I__4040 (
            .O(N__20289),
            .I(\Lab_UT.dictrl.N_5 ));
    InMux I__4039 (
            .O(N__20284),
            .I(N__20280));
    InMux I__4038 (
            .O(N__20283),
            .I(N__20277));
    LocalMux I__4037 (
            .O(N__20280),
            .I(N__20274));
    LocalMux I__4036 (
            .O(N__20277),
            .I(N__20271));
    Span4Mux_h I__4035 (
            .O(N__20274),
            .I(N__20268));
    Odrv4 I__4034 (
            .O(N__20271),
            .I(\Lab_UT.dictrl.N_6 ));
    Odrv4 I__4033 (
            .O(N__20268),
            .I(\Lab_UT.dictrl.N_6 ));
    CascadeMux I__4032 (
            .O(N__20263),
            .I(\Lab_UT.dictrl.r_enable2_3_iv_0_cascade_ ));
    InMux I__4031 (
            .O(N__20260),
            .I(N__20257));
    LocalMux I__4030 (
            .O(N__20257),
            .I(N__20254));
    Odrv4 I__4029 (
            .O(N__20254),
            .I(\Lab_UT.dictrl.r_enable2_3_iv_3 ));
    InMux I__4028 (
            .O(N__20251),
            .I(N__20248));
    LocalMux I__4027 (
            .O(N__20248),
            .I(N__20245));
    Span4Mux_h I__4026 (
            .O(N__20245),
            .I(N__20242));
    Sp12to4 I__4025 (
            .O(N__20242),
            .I(N__20239));
    Odrv12 I__4024 (
            .O(N__20239),
            .I(\Lab_UT.dictrl.r_Sone_init17_4 ));
    InMux I__4023 (
            .O(N__20236),
            .I(N__20230));
    InMux I__4022 (
            .O(N__20235),
            .I(N__20230));
    LocalMux I__4021 (
            .O(N__20230),
            .I(\Lab_UT.dictrl.r_dicLdMtens23_i_6 ));
    CascadeMux I__4020 (
            .O(N__20227),
            .I(\Lab_UT.dictrl.un1_r_dicLdMtens19_0_cascade_ ));
    InMux I__4019 (
            .O(N__20224),
            .I(N__20220));
    InMux I__4018 (
            .O(N__20223),
            .I(N__20217));
    LocalMux I__4017 (
            .O(N__20220),
            .I(\Lab_UT.dictrl.r_alarm_or_timeZ0 ));
    LocalMux I__4016 (
            .O(N__20217),
            .I(\Lab_UT.dictrl.r_alarm_or_timeZ0 ));
    InMux I__4015 (
            .O(N__20212),
            .I(N__20209));
    LocalMux I__4014 (
            .O(N__20209),
            .I(\Lab_UT.dictrl.r_dicLdMtens18_i_6 ));
    InMux I__4013 (
            .O(N__20206),
            .I(N__20203));
    LocalMux I__4012 (
            .O(N__20203),
            .I(\Lab_UT.dictrl.r_dicLdMtens17_i_6 ));
    InMux I__4011 (
            .O(N__20200),
            .I(N__20197));
    LocalMux I__4010 (
            .O(N__20197),
            .I(N__20194));
    Odrv4 I__4009 (
            .O(N__20194),
            .I(\Lab_UT.dictrl.r_enable1_2_m ));
    CascadeMux I__4008 (
            .O(N__20191),
            .I(\Lab_UT.dictrl.r_enable1_2_m_cascade_ ));
    InMux I__4007 (
            .O(N__20188),
            .I(N__20185));
    LocalMux I__4006 (
            .O(N__20185),
            .I(N__20182));
    Odrv12 I__4005 (
            .O(N__20182),
            .I(\Lab_UT.dictrl.g0_i_a4_0 ));
    InMux I__4004 (
            .O(N__20179),
            .I(N__20173));
    InMux I__4003 (
            .O(N__20178),
            .I(N__20173));
    LocalMux I__4002 (
            .O(N__20173),
            .I(\Lab_UT.dictrl.r_enableZ0Z2 ));
    InMux I__4001 (
            .O(N__20170),
            .I(N__20161));
    InMux I__4000 (
            .O(N__20169),
            .I(N__20154));
    InMux I__3999 (
            .O(N__20168),
            .I(N__20154));
    InMux I__3998 (
            .O(N__20167),
            .I(N__20154));
    InMux I__3997 (
            .O(N__20166),
            .I(N__20147));
    InMux I__3996 (
            .O(N__20165),
            .I(N__20147));
    InMux I__3995 (
            .O(N__20164),
            .I(N__20147));
    LocalMux I__3994 (
            .O(N__20161),
            .I(N__20144));
    LocalMux I__3993 (
            .O(N__20154),
            .I(N__20141));
    LocalMux I__3992 (
            .O(N__20147),
            .I(N__20138));
    Span4Mux_v I__3991 (
            .O(N__20144),
            .I(N__20135));
    Span4Mux_v I__3990 (
            .O(N__20141),
            .I(N__20130));
    Span4Mux_h I__3989 (
            .O(N__20138),
            .I(N__20130));
    Odrv4 I__3988 (
            .O(N__20135),
            .I(\Lab_UT.dictrl.enableSeg2 ));
    Odrv4 I__3987 (
            .O(N__20130),
            .I(\Lab_UT.dictrl.enableSeg2 ));
    InMux I__3986 (
            .O(N__20125),
            .I(N__20122));
    LocalMux I__3985 (
            .O(N__20122),
            .I(\Lab_UT.dictrl.currState_0_ret_20and_1_0 ));
    InMux I__3984 (
            .O(N__20119),
            .I(N__20115));
    InMux I__3983 (
            .O(N__20118),
            .I(N__20112));
    LocalMux I__3982 (
            .O(N__20115),
            .I(\Lab_UT.dictrl.r_dicLdMtens16_reti ));
    LocalMux I__3981 (
            .O(N__20112),
            .I(\Lab_UT.dictrl.r_dicLdMtens16_reti ));
    InMux I__3980 (
            .O(N__20107),
            .I(N__20103));
    InMux I__3979 (
            .O(N__20106),
            .I(N__20100));
    LocalMux I__3978 (
            .O(N__20103),
            .I(N__20095));
    LocalMux I__3977 (
            .O(N__20100),
            .I(N__20095));
    Span4Mux_v I__3976 (
            .O(N__20095),
            .I(N__20092));
    Span4Mux_h I__3975 (
            .O(N__20092),
            .I(N__20089));
    Odrv4 I__3974 (
            .O(N__20089),
            .I(\Lab_UT.dictrl.r_dicLdMtens19 ));
    InMux I__3973 (
            .O(N__20086),
            .I(N__20083));
    LocalMux I__3972 (
            .O(N__20083),
            .I(N__20080));
    Odrv12 I__3971 (
            .O(N__20080),
            .I(\Lab_UT.dictrl.r_dicLdMtens22_i_6 ));
    InMux I__3970 (
            .O(N__20077),
            .I(N__20062));
    InMux I__3969 (
            .O(N__20076),
            .I(N__20062));
    InMux I__3968 (
            .O(N__20075),
            .I(N__20062));
    InMux I__3967 (
            .O(N__20074),
            .I(N__20062));
    InMux I__3966 (
            .O(N__20073),
            .I(N__20055));
    InMux I__3965 (
            .O(N__20072),
            .I(N__20055));
    InMux I__3964 (
            .O(N__20071),
            .I(N__20055));
    LocalMux I__3963 (
            .O(N__20062),
            .I(N__20052));
    LocalMux I__3962 (
            .O(N__20055),
            .I(\Lab_UT.Sten_at_1 ));
    Odrv4 I__3961 (
            .O(N__20052),
            .I(\Lab_UT.Sten_at_1 ));
    InMux I__3960 (
            .O(N__20047),
            .I(N__20031));
    InMux I__3959 (
            .O(N__20046),
            .I(N__20031));
    InMux I__3958 (
            .O(N__20045),
            .I(N__20031));
    InMux I__3957 (
            .O(N__20044),
            .I(N__20031));
    InMux I__3956 (
            .O(N__20043),
            .I(N__20021));
    InMux I__3955 (
            .O(N__20042),
            .I(N__20021));
    InMux I__3954 (
            .O(N__20041),
            .I(N__20021));
    InMux I__3953 (
            .O(N__20040),
            .I(N__20021));
    LocalMux I__3952 (
            .O(N__20031),
            .I(N__20018));
    InMux I__3951 (
            .O(N__20030),
            .I(N__20015));
    LocalMux I__3950 (
            .O(N__20021),
            .I(\Lab_UT.Sten_at_0 ));
    Odrv4 I__3949 (
            .O(N__20018),
            .I(\Lab_UT.Sten_at_0 ));
    LocalMux I__3948 (
            .O(N__20015),
            .I(\Lab_UT.Sten_at_0 ));
    CascadeMux I__3947 (
            .O(N__20008),
            .I(N__20002));
    InMux I__3946 (
            .O(N__20007),
            .I(N__19993));
    InMux I__3945 (
            .O(N__20006),
            .I(N__19993));
    InMux I__3944 (
            .O(N__20005),
            .I(N__19993));
    InMux I__3943 (
            .O(N__20002),
            .I(N__19993));
    LocalMux I__3942 (
            .O(N__19993),
            .I(N__19988));
    CascadeMux I__3941 (
            .O(N__19992),
            .I(N__19984));
    CascadeMux I__3940 (
            .O(N__19991),
            .I(N__19980));
    Span4Mux_h I__3939 (
            .O(N__19988),
            .I(N__19976));
    InMux I__3938 (
            .O(N__19987),
            .I(N__19973));
    InMux I__3937 (
            .O(N__19984),
            .I(N__19966));
    InMux I__3936 (
            .O(N__19983),
            .I(N__19966));
    InMux I__3935 (
            .O(N__19980),
            .I(N__19966));
    InMux I__3934 (
            .O(N__19979),
            .I(N__19963));
    Odrv4 I__3933 (
            .O(N__19976),
            .I(\Lab_UT.Sten_at_3 ));
    LocalMux I__3932 (
            .O(N__19973),
            .I(\Lab_UT.Sten_at_3 ));
    LocalMux I__3931 (
            .O(N__19966),
            .I(\Lab_UT.Sten_at_3 ));
    LocalMux I__3930 (
            .O(N__19963),
            .I(\Lab_UT.Sten_at_3 ));
    CascadeMux I__3929 (
            .O(N__19954),
            .I(\Lab_UT.Sten_at_1_cascade_ ));
    CascadeMux I__3928 (
            .O(N__19951),
            .I(N__19945));
    CascadeMux I__3927 (
            .O(N__19950),
            .I(N__19942));
    CascadeMux I__3926 (
            .O(N__19949),
            .I(N__19939));
    CascadeMux I__3925 (
            .O(N__19948),
            .I(N__19934));
    InMux I__3924 (
            .O(N__19945),
            .I(N__19924));
    InMux I__3923 (
            .O(N__19942),
            .I(N__19924));
    InMux I__3922 (
            .O(N__19939),
            .I(N__19924));
    InMux I__3921 (
            .O(N__19938),
            .I(N__19924));
    InMux I__3920 (
            .O(N__19937),
            .I(N__19916));
    InMux I__3919 (
            .O(N__19934),
            .I(N__19916));
    InMux I__3918 (
            .O(N__19933),
            .I(N__19916));
    LocalMux I__3917 (
            .O(N__19924),
            .I(N__19913));
    InMux I__3916 (
            .O(N__19923),
            .I(N__19910));
    LocalMux I__3915 (
            .O(N__19916),
            .I(\Lab_UT.Sten_at_2 ));
    Odrv4 I__3914 (
            .O(N__19913),
            .I(\Lab_UT.Sten_at_2 ));
    LocalMux I__3913 (
            .O(N__19910),
            .I(\Lab_UT.Sten_at_2 ));
    InMux I__3912 (
            .O(N__19903),
            .I(N__19900));
    LocalMux I__3911 (
            .O(N__19900),
            .I(\Lab_UT.segmentUQ_0_0_0 ));
    CascadeMux I__3910 (
            .O(N__19897),
            .I(N__19890));
    InMux I__3909 (
            .O(N__19896),
            .I(N__19870));
    InMux I__3908 (
            .O(N__19895),
            .I(N__19870));
    InMux I__3907 (
            .O(N__19894),
            .I(N__19865));
    InMux I__3906 (
            .O(N__19893),
            .I(N__19865));
    InMux I__3905 (
            .O(N__19890),
            .I(N__19858));
    InMux I__3904 (
            .O(N__19889),
            .I(N__19858));
    InMux I__3903 (
            .O(N__19888),
            .I(N__19858));
    CascadeMux I__3902 (
            .O(N__19887),
            .I(N__19852));
    InMux I__3901 (
            .O(N__19886),
            .I(N__19845));
    InMux I__3900 (
            .O(N__19885),
            .I(N__19840));
    InMux I__3899 (
            .O(N__19884),
            .I(N__19840));
    InMux I__3898 (
            .O(N__19883),
            .I(N__19835));
    InMux I__3897 (
            .O(N__19882),
            .I(N__19835));
    InMux I__3896 (
            .O(N__19881),
            .I(N__19828));
    InMux I__3895 (
            .O(N__19880),
            .I(N__19828));
    InMux I__3894 (
            .O(N__19879),
            .I(N__19828));
    InMux I__3893 (
            .O(N__19878),
            .I(N__19821));
    InMux I__3892 (
            .O(N__19877),
            .I(N__19821));
    InMux I__3891 (
            .O(N__19876),
            .I(N__19821));
    CascadeMux I__3890 (
            .O(N__19875),
            .I(N__19817));
    LocalMux I__3889 (
            .O(N__19870),
            .I(N__19810));
    LocalMux I__3888 (
            .O(N__19865),
            .I(N__19810));
    LocalMux I__3887 (
            .O(N__19858),
            .I(N__19810));
    InMux I__3886 (
            .O(N__19857),
            .I(N__19807));
    InMux I__3885 (
            .O(N__19856),
            .I(N__19802));
    InMux I__3884 (
            .O(N__19855),
            .I(N__19802));
    InMux I__3883 (
            .O(N__19852),
            .I(N__19797));
    InMux I__3882 (
            .O(N__19851),
            .I(N__19797));
    InMux I__3881 (
            .O(N__19850),
            .I(N__19790));
    InMux I__3880 (
            .O(N__19849),
            .I(N__19790));
    InMux I__3879 (
            .O(N__19848),
            .I(N__19790));
    LocalMux I__3878 (
            .O(N__19845),
            .I(N__19783));
    LocalMux I__3877 (
            .O(N__19840),
            .I(N__19783));
    LocalMux I__3876 (
            .O(N__19835),
            .I(N__19783));
    LocalMux I__3875 (
            .O(N__19828),
            .I(N__19778));
    LocalMux I__3874 (
            .O(N__19821),
            .I(N__19778));
    InMux I__3873 (
            .O(N__19820),
            .I(N__19773));
    InMux I__3872 (
            .O(N__19817),
            .I(N__19773));
    Span4Mux_v I__3871 (
            .O(N__19810),
            .I(N__19770));
    LocalMux I__3870 (
            .O(N__19807),
            .I(N__19761));
    LocalMux I__3869 (
            .O(N__19802),
            .I(N__19761));
    LocalMux I__3868 (
            .O(N__19797),
            .I(N__19761));
    LocalMux I__3867 (
            .O(N__19790),
            .I(N__19761));
    Span4Mux_h I__3866 (
            .O(N__19783),
            .I(N__19758));
    Span4Mux_h I__3865 (
            .O(N__19778),
            .I(N__19755));
    LocalMux I__3864 (
            .O(N__19773),
            .I(N__19750));
    Span4Mux_h I__3863 (
            .O(N__19770),
            .I(N__19750));
    Odrv4 I__3862 (
            .O(N__19761),
            .I(\Lab_UT.dictrl.L3_segment1_1 ));
    Odrv4 I__3861 (
            .O(N__19758),
            .I(\Lab_UT.dictrl.L3_segment1_1 ));
    Odrv4 I__3860 (
            .O(N__19755),
            .I(\Lab_UT.dictrl.L3_segment1_1 ));
    Odrv4 I__3859 (
            .O(N__19750),
            .I(\Lab_UT.dictrl.L3_segment1_1 ));
    CascadeMux I__3858 (
            .O(N__19741),
            .I(N__19733));
    CascadeMux I__3857 (
            .O(N__19740),
            .I(N__19730));
    CascadeMux I__3856 (
            .O(N__19739),
            .I(N__19727));
    CascadeMux I__3855 (
            .O(N__19738),
            .I(N__19723));
    InMux I__3854 (
            .O(N__19737),
            .I(N__19713));
    InMux I__3853 (
            .O(N__19736),
            .I(N__19713));
    InMux I__3852 (
            .O(N__19733),
            .I(N__19713));
    InMux I__3851 (
            .O(N__19730),
            .I(N__19713));
    InMux I__3850 (
            .O(N__19727),
            .I(N__19704));
    InMux I__3849 (
            .O(N__19726),
            .I(N__19704));
    InMux I__3848 (
            .O(N__19723),
            .I(N__19704));
    InMux I__3847 (
            .O(N__19722),
            .I(N__19704));
    LocalMux I__3846 (
            .O(N__19713),
            .I(N__19699));
    LocalMux I__3845 (
            .O(N__19704),
            .I(N__19699));
    Odrv4 I__3844 (
            .O(N__19699),
            .I(\Lab_UT.Sone_at_1 ));
    InMux I__3843 (
            .O(N__19696),
            .I(N__19690));
    InMux I__3842 (
            .O(N__19695),
            .I(N__19690));
    LocalMux I__3841 (
            .O(N__19690),
            .I(N__19687));
    Odrv4 I__3840 (
            .O(N__19687),
            .I(\Lab_UT.dictrl.r_enable1_2_i_m ));
    InMux I__3839 (
            .O(N__19684),
            .I(N__19672));
    InMux I__3838 (
            .O(N__19683),
            .I(N__19672));
    InMux I__3837 (
            .O(N__19682),
            .I(N__19672));
    InMux I__3836 (
            .O(N__19681),
            .I(N__19672));
    LocalMux I__3835 (
            .O(N__19672),
            .I(N__19661));
    InMux I__3834 (
            .O(N__19671),
            .I(N__19646));
    InMux I__3833 (
            .O(N__19670),
            .I(N__19646));
    InMux I__3832 (
            .O(N__19669),
            .I(N__19646));
    InMux I__3831 (
            .O(N__19668),
            .I(N__19646));
    InMux I__3830 (
            .O(N__19667),
            .I(N__19646));
    InMux I__3829 (
            .O(N__19666),
            .I(N__19646));
    InMux I__3828 (
            .O(N__19665),
            .I(N__19639));
    InMux I__3827 (
            .O(N__19664),
            .I(N__19639));
    Span4Mux_v I__3826 (
            .O(N__19661),
            .I(N__19636));
    InMux I__3825 (
            .O(N__19660),
            .I(N__19631));
    InMux I__3824 (
            .O(N__19659),
            .I(N__19631));
    LocalMux I__3823 (
            .O(N__19646),
            .I(N__19628));
    InMux I__3822 (
            .O(N__19645),
            .I(N__19623));
    InMux I__3821 (
            .O(N__19644),
            .I(N__19623));
    LocalMux I__3820 (
            .O(N__19639),
            .I(\Lab_UT.alarm_or_time_0 ));
    Odrv4 I__3819 (
            .O(N__19636),
            .I(\Lab_UT.alarm_or_time_0 ));
    LocalMux I__3818 (
            .O(N__19631),
            .I(\Lab_UT.alarm_or_time_0 ));
    Odrv4 I__3817 (
            .O(N__19628),
            .I(\Lab_UT.alarm_or_time_0 ));
    LocalMux I__3816 (
            .O(N__19623),
            .I(\Lab_UT.alarm_or_time_0 ));
    CascadeMux I__3815 (
            .O(N__19612),
            .I(\Lab_UT.alarm_or_time_0_cascade_ ));
    CascadeMux I__3814 (
            .O(N__19609),
            .I(N__19605));
    InMux I__3813 (
            .O(N__19608),
            .I(N__19594));
    InMux I__3812 (
            .O(N__19605),
            .I(N__19594));
    InMux I__3811 (
            .O(N__19604),
            .I(N__19594));
    InMux I__3810 (
            .O(N__19603),
            .I(N__19594));
    LocalMux I__3809 (
            .O(N__19594),
            .I(N__19591));
    Span4Mux_h I__3808 (
            .O(N__19591),
            .I(N__19584));
    InMux I__3807 (
            .O(N__19590),
            .I(N__19581));
    InMux I__3806 (
            .O(N__19589),
            .I(N__19576));
    InMux I__3805 (
            .O(N__19588),
            .I(N__19576));
    InMux I__3804 (
            .O(N__19587),
            .I(N__19573));
    Odrv4 I__3803 (
            .O(N__19584),
            .I(\Lab_UT.Mten_at_2 ));
    LocalMux I__3802 (
            .O(N__19581),
            .I(\Lab_UT.Mten_at_2 ));
    LocalMux I__3801 (
            .O(N__19576),
            .I(\Lab_UT.Mten_at_2 ));
    LocalMux I__3800 (
            .O(N__19573),
            .I(\Lab_UT.Mten_at_2 ));
    InMux I__3799 (
            .O(N__19564),
            .I(N__19556));
    InMux I__3798 (
            .O(N__19563),
            .I(N__19549));
    InMux I__3797 (
            .O(N__19562),
            .I(N__19549));
    InMux I__3796 (
            .O(N__19561),
            .I(N__19549));
    InMux I__3795 (
            .O(N__19560),
            .I(N__19544));
    InMux I__3794 (
            .O(N__19559),
            .I(N__19544));
    LocalMux I__3793 (
            .O(N__19556),
            .I(N__19536));
    LocalMux I__3792 (
            .O(N__19549),
            .I(N__19536));
    LocalMux I__3791 (
            .O(N__19544),
            .I(N__19536));
    InMux I__3790 (
            .O(N__19543),
            .I(N__19533));
    Span4Mux_h I__3789 (
            .O(N__19536),
            .I(N__19530));
    LocalMux I__3788 (
            .O(N__19533),
            .I(N__19527));
    Odrv4 I__3787 (
            .O(N__19530),
            .I(\Lab_UT.dictrl.enableSeg1 ));
    Odrv12 I__3786 (
            .O(N__19527),
            .I(\Lab_UT.dictrl.enableSeg1 ));
    CascadeMux I__3785 (
            .O(N__19522),
            .I(\Lab_UT.L3_segment1_1_2_cascade_ ));
    InMux I__3784 (
            .O(N__19519),
            .I(N__19516));
    LocalMux I__3783 (
            .O(N__19516),
            .I(\uu2.bitmapZ0Z_93 ));
    InMux I__3782 (
            .O(N__19513),
            .I(N__19510));
    LocalMux I__3781 (
            .O(N__19510),
            .I(\uu2.bitmap_pmux_25_bm_1 ));
    CascadeMux I__3780 (
            .O(N__19507),
            .I(N__19504));
    InMux I__3779 (
            .O(N__19504),
            .I(N__19501));
    LocalMux I__3778 (
            .O(N__19501),
            .I(\uu2.bitmapZ0Z_221 ));
    CascadeMux I__3777 (
            .O(N__19498),
            .I(N__19488));
    CascadeMux I__3776 (
            .O(N__19497),
            .I(N__19484));
    InMux I__3775 (
            .O(N__19496),
            .I(N__19480));
    InMux I__3774 (
            .O(N__19495),
            .I(N__19477));
    InMux I__3773 (
            .O(N__19494),
            .I(N__19474));
    InMux I__3772 (
            .O(N__19493),
            .I(N__19468));
    InMux I__3771 (
            .O(N__19492),
            .I(N__19468));
    InMux I__3770 (
            .O(N__19491),
            .I(N__19465));
    InMux I__3769 (
            .O(N__19488),
            .I(N__19460));
    InMux I__3768 (
            .O(N__19487),
            .I(N__19460));
    InMux I__3767 (
            .O(N__19484),
            .I(N__19453));
    InMux I__3766 (
            .O(N__19483),
            .I(N__19453));
    LocalMux I__3765 (
            .O(N__19480),
            .I(N__19448));
    LocalMux I__3764 (
            .O(N__19477),
            .I(N__19448));
    LocalMux I__3763 (
            .O(N__19474),
            .I(N__19445));
    InMux I__3762 (
            .O(N__19473),
            .I(N__19442));
    LocalMux I__3761 (
            .O(N__19468),
            .I(N__19439));
    LocalMux I__3760 (
            .O(N__19465),
            .I(N__19432));
    LocalMux I__3759 (
            .O(N__19460),
            .I(N__19429));
    CascadeMux I__3758 (
            .O(N__19459),
            .I(N__19426));
    CascadeMux I__3757 (
            .O(N__19458),
            .I(N__19422));
    LocalMux I__3756 (
            .O(N__19453),
            .I(N__19415));
    Span4Mux_h I__3755 (
            .O(N__19448),
            .I(N__19415));
    Span4Mux_h I__3754 (
            .O(N__19445),
            .I(N__19415));
    LocalMux I__3753 (
            .O(N__19442),
            .I(N__19410));
    Span4Mux_h I__3752 (
            .O(N__19439),
            .I(N__19410));
    InMux I__3751 (
            .O(N__19438),
            .I(N__19407));
    InMux I__3750 (
            .O(N__19437),
            .I(N__19402));
    InMux I__3749 (
            .O(N__19436),
            .I(N__19402));
    InMux I__3748 (
            .O(N__19435),
            .I(N__19399));
    Span4Mux_h I__3747 (
            .O(N__19432),
            .I(N__19394));
    Span4Mux_h I__3746 (
            .O(N__19429),
            .I(N__19394));
    InMux I__3745 (
            .O(N__19426),
            .I(N__19391));
    InMux I__3744 (
            .O(N__19425),
            .I(N__19386));
    InMux I__3743 (
            .O(N__19422),
            .I(N__19386));
    Odrv4 I__3742 (
            .O(N__19415),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    Odrv4 I__3741 (
            .O(N__19410),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    LocalMux I__3740 (
            .O(N__19407),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    LocalMux I__3739 (
            .O(N__19402),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    LocalMux I__3738 (
            .O(N__19399),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    Odrv4 I__3737 (
            .O(N__19394),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    LocalMux I__3736 (
            .O(N__19391),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    LocalMux I__3735 (
            .O(N__19386),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    InMux I__3734 (
            .O(N__19369),
            .I(N__19366));
    LocalMux I__3733 (
            .O(N__19366),
            .I(N__19363));
    Odrv4 I__3732 (
            .O(N__19363),
            .I(\uu2.bitmap_RNI1D952Z0Z_93 ));
    InMux I__3731 (
            .O(N__19360),
            .I(N__19344));
    InMux I__3730 (
            .O(N__19359),
            .I(N__19344));
    InMux I__3729 (
            .O(N__19358),
            .I(N__19344));
    InMux I__3728 (
            .O(N__19357),
            .I(N__19344));
    InMux I__3727 (
            .O(N__19356),
            .I(N__19335));
    InMux I__3726 (
            .O(N__19355),
            .I(N__19335));
    InMux I__3725 (
            .O(N__19354),
            .I(N__19335));
    InMux I__3724 (
            .O(N__19353),
            .I(N__19335));
    LocalMux I__3723 (
            .O(N__19344),
            .I(\Lab_UT.Sone_at_0 ));
    LocalMux I__3722 (
            .O(N__19335),
            .I(\Lab_UT.Sone_at_0 ));
    CascadeMux I__3721 (
            .O(N__19330),
            .I(\Lab_UT.Sone_at_0_cascade_ ));
    InMux I__3720 (
            .O(N__19327),
            .I(N__19324));
    LocalMux I__3719 (
            .O(N__19324),
            .I(N__19321));
    Odrv4 I__3718 (
            .O(N__19321),
            .I(\Lab_UT.N_77_2 ));
    CascadeMux I__3717 (
            .O(N__19318),
            .I(N__19312));
    CascadeMux I__3716 (
            .O(N__19317),
            .I(N__19307));
    CascadeMux I__3715 (
            .O(N__19316),
            .I(N__19301));
    CascadeMux I__3714 (
            .O(N__19315),
            .I(N__19298));
    InMux I__3713 (
            .O(N__19312),
            .I(N__19289));
    InMux I__3712 (
            .O(N__19311),
            .I(N__19289));
    InMux I__3711 (
            .O(N__19310),
            .I(N__19289));
    InMux I__3710 (
            .O(N__19307),
            .I(N__19289));
    InMux I__3709 (
            .O(N__19306),
            .I(N__19286));
    InMux I__3708 (
            .O(N__19305),
            .I(N__19277));
    InMux I__3707 (
            .O(N__19304),
            .I(N__19277));
    InMux I__3706 (
            .O(N__19301),
            .I(N__19277));
    InMux I__3705 (
            .O(N__19298),
            .I(N__19277));
    LocalMux I__3704 (
            .O(N__19289),
            .I(\Lab_UT.Sone_at_3 ));
    LocalMux I__3703 (
            .O(N__19286),
            .I(\Lab_UT.Sone_at_3 ));
    LocalMux I__3702 (
            .O(N__19277),
            .I(\Lab_UT.Sone_at_3 ));
    InMux I__3701 (
            .O(N__19270),
            .I(N__19254));
    InMux I__3700 (
            .O(N__19269),
            .I(N__19254));
    InMux I__3699 (
            .O(N__19268),
            .I(N__19254));
    InMux I__3698 (
            .O(N__19267),
            .I(N__19254));
    InMux I__3697 (
            .O(N__19266),
            .I(N__19245));
    InMux I__3696 (
            .O(N__19265),
            .I(N__19245));
    InMux I__3695 (
            .O(N__19264),
            .I(N__19245));
    InMux I__3694 (
            .O(N__19263),
            .I(N__19245));
    LocalMux I__3693 (
            .O(N__19254),
            .I(\Lab_UT.Sone_at_2 ));
    LocalMux I__3692 (
            .O(N__19245),
            .I(\Lab_UT.Sone_at_2 ));
    InMux I__3691 (
            .O(N__19240),
            .I(N__19231));
    InMux I__3690 (
            .O(N__19239),
            .I(N__19231));
    InMux I__3689 (
            .O(N__19238),
            .I(N__19231));
    LocalMux I__3688 (
            .O(N__19231),
            .I(\resetGen.reset_countZ0Z_1 ));
    InMux I__3687 (
            .O(N__19228),
            .I(N__19219));
    InMux I__3686 (
            .O(N__19227),
            .I(N__19219));
    InMux I__3685 (
            .O(N__19226),
            .I(N__19219));
    LocalMux I__3684 (
            .O(N__19219),
            .I(N__19215));
    InMux I__3683 (
            .O(N__19218),
            .I(N__19212));
    Span4Mux_h I__3682 (
            .O(N__19215),
            .I(N__19209));
    LocalMux I__3681 (
            .O(N__19212),
            .I(\resetGen.reset_countZ0Z_0 ));
    Odrv4 I__3680 (
            .O(N__19209),
            .I(\resetGen.reset_countZ0Z_0 ));
    InMux I__3679 (
            .O(N__19204),
            .I(N__19201));
    LocalMux I__3678 (
            .O(N__19201),
            .I(N__19198));
    Span4Mux_h I__3677 (
            .O(N__19198),
            .I(N__19195));
    Odrv4 I__3676 (
            .O(N__19195),
            .I(\resetGen.un241_ci ));
    CascadeMux I__3675 (
            .O(N__19192),
            .I(N__19188));
    InMux I__3674 (
            .O(N__19191),
            .I(N__19183));
    InMux I__3673 (
            .O(N__19188),
            .I(N__19176));
    InMux I__3672 (
            .O(N__19187),
            .I(N__19176));
    InMux I__3671 (
            .O(N__19186),
            .I(N__19176));
    LocalMux I__3670 (
            .O(N__19183),
            .I(N__19173));
    LocalMux I__3669 (
            .O(N__19176),
            .I(N__19168));
    Span4Mux_v I__3668 (
            .O(N__19173),
            .I(N__19165));
    InMux I__3667 (
            .O(N__19172),
            .I(N__19162));
    InMux I__3666 (
            .O(N__19171),
            .I(N__19159));
    Span4Mux_v I__3665 (
            .O(N__19168),
            .I(N__19154));
    Span4Mux_v I__3664 (
            .O(N__19165),
            .I(N__19154));
    LocalMux I__3663 (
            .O(N__19162),
            .I(\resetGen.reset_countZ0Z_4 ));
    LocalMux I__3662 (
            .O(N__19159),
            .I(\resetGen.reset_countZ0Z_4 ));
    Odrv4 I__3661 (
            .O(N__19154),
            .I(\resetGen.reset_countZ0Z_4 ));
    CascadeMux I__3660 (
            .O(N__19147),
            .I(\resetGen.un241_ci_cascade_ ));
    InMux I__3659 (
            .O(N__19144),
            .I(N__19141));
    LocalMux I__3658 (
            .O(N__19141),
            .I(N__19136));
    InMux I__3657 (
            .O(N__19140),
            .I(N__19131));
    InMux I__3656 (
            .O(N__19139),
            .I(N__19131));
    Span4Mux_h I__3655 (
            .O(N__19136),
            .I(N__19128));
    LocalMux I__3654 (
            .O(N__19131),
            .I(\resetGen.reset_countZ0Z_2 ));
    Odrv4 I__3653 (
            .O(N__19128),
            .I(\resetGen.reset_countZ0Z_2 ));
    InMux I__3652 (
            .O(N__19123),
            .I(N__19120));
    LocalMux I__3651 (
            .O(N__19120),
            .I(N__19117));
    Span4Mux_v I__3650 (
            .O(N__19117),
            .I(N__19114));
    Odrv4 I__3649 (
            .O(N__19114),
            .I(\Lab_UT.uu0.delay_lineZ0Z_1 ));
    IoInMux I__3648 (
            .O(N__19111),
            .I(N__19108));
    LocalMux I__3647 (
            .O(N__19108),
            .I(N__19105));
    Span4Mux_s0_h I__3646 (
            .O(N__19105),
            .I(N__19102));
    Span4Mux_h I__3645 (
            .O(N__19102),
            .I(N__19099));
    Odrv4 I__3644 (
            .O(N__19099),
            .I(\Lab_UT.uu0.un11_l_count_i ));
    InMux I__3643 (
            .O(N__19096),
            .I(N__19093));
    LocalMux I__3642 (
            .O(N__19093),
            .I(N__19090));
    Odrv4 I__3641 (
            .O(N__19090),
            .I(\Lab_UT.L3_segment1_1_0_3 ));
    CascadeMux I__3640 (
            .O(N__19087),
            .I(\Lab_UT.L3_segment1_0_i_1_0_cascade_ ));
    InMux I__3639 (
            .O(N__19084),
            .I(N__19081));
    LocalMux I__3638 (
            .O(N__19081),
            .I(N__19078));
    Odrv12 I__3637 (
            .O(N__19078),
            .I(\uu2.bitmapZ0Z_58 ));
    InMux I__3636 (
            .O(N__19075),
            .I(N__19072));
    LocalMux I__3635 (
            .O(N__19072),
            .I(\Lab_UT.L3_segment1_0_i_1_1 ));
    CascadeMux I__3634 (
            .O(N__19069),
            .I(N__19065));
    InMux I__3633 (
            .O(N__19068),
            .I(N__19051));
    InMux I__3632 (
            .O(N__19065),
            .I(N__19051));
    InMux I__3631 (
            .O(N__19064),
            .I(N__19051));
    InMux I__3630 (
            .O(N__19063),
            .I(N__19051));
    InMux I__3629 (
            .O(N__19062),
            .I(N__19051));
    LocalMux I__3628 (
            .O(N__19051),
            .I(N__19046));
    InMux I__3627 (
            .O(N__19050),
            .I(N__19041));
    InMux I__3626 (
            .O(N__19049),
            .I(N__19041));
    Odrv4 I__3625 (
            .O(N__19046),
            .I(\uu2.w_addr_userZ0Z_0 ));
    LocalMux I__3624 (
            .O(N__19041),
            .I(\uu2.w_addr_userZ0Z_0 ));
    CascadeMux I__3623 (
            .O(N__19036),
            .I(N__19031));
    InMux I__3622 (
            .O(N__19035),
            .I(N__19027));
    CascadeMux I__3621 (
            .O(N__19034),
            .I(N__19024));
    InMux I__3620 (
            .O(N__19031),
            .I(N__19018));
    InMux I__3619 (
            .O(N__19030),
            .I(N__19018));
    LocalMux I__3618 (
            .O(N__19027),
            .I(N__19015));
    InMux I__3617 (
            .O(N__19024),
            .I(N__19010));
    InMux I__3616 (
            .O(N__19023),
            .I(N__19010));
    LocalMux I__3615 (
            .O(N__19018),
            .I(N__19007));
    Span4Mux_s3_v I__3614 (
            .O(N__19015),
            .I(N__19004));
    LocalMux I__3613 (
            .O(N__19010),
            .I(\uu2.w_addr_userZ0Z_2 ));
    Odrv4 I__3612 (
            .O(N__19007),
            .I(\uu2.w_addr_userZ0Z_2 ));
    Odrv4 I__3611 (
            .O(N__19004),
            .I(\uu2.w_addr_userZ0Z_2 ));
    CascadeMux I__3610 (
            .O(N__18997),
            .I(N__18994));
    InMux I__3609 (
            .O(N__18994),
            .I(N__18988));
    InMux I__3608 (
            .O(N__18993),
            .I(N__18983));
    InMux I__3607 (
            .O(N__18992),
            .I(N__18983));
    InMux I__3606 (
            .O(N__18991),
            .I(N__18980));
    LocalMux I__3605 (
            .O(N__18988),
            .I(\uu2.w_addr_userZ0Z_3 ));
    LocalMux I__3604 (
            .O(N__18983),
            .I(\uu2.w_addr_userZ0Z_3 ));
    LocalMux I__3603 (
            .O(N__18980),
            .I(\uu2.w_addr_userZ0Z_3 ));
    InMux I__3602 (
            .O(N__18973),
            .I(N__18970));
    LocalMux I__3601 (
            .O(N__18970),
            .I(N__18964));
    InMux I__3600 (
            .O(N__18969),
            .I(N__18955));
    InMux I__3599 (
            .O(N__18968),
            .I(N__18955));
    InMux I__3598 (
            .O(N__18967),
            .I(N__18955));
    Span4Mux_h I__3597 (
            .O(N__18964),
            .I(N__18952));
    InMux I__3596 (
            .O(N__18963),
            .I(N__18947));
    InMux I__3595 (
            .O(N__18962),
            .I(N__18947));
    LocalMux I__3594 (
            .O(N__18955),
            .I(\uu2.w_addr_userZ0Z_1 ));
    Odrv4 I__3593 (
            .O(N__18952),
            .I(\uu2.w_addr_userZ0Z_1 ));
    LocalMux I__3592 (
            .O(N__18947),
            .I(\uu2.w_addr_userZ0Z_1 ));
    CascadeMux I__3591 (
            .O(N__18940),
            .I(\resetGen.un252_ci_cascade_ ));
    InMux I__3590 (
            .O(N__18937),
            .I(N__18934));
    LocalMux I__3589 (
            .O(N__18934),
            .I(N__18930));
    InMux I__3588 (
            .O(N__18933),
            .I(N__18927));
    Span4Mux_v I__3587 (
            .O(N__18930),
            .I(N__18924));
    LocalMux I__3586 (
            .O(N__18927),
            .I(\resetGen.reset_countZ0Z_3 ));
    Odrv4 I__3585 (
            .O(N__18924),
            .I(\resetGen.reset_countZ0Z_3 ));
    CEMux I__3584 (
            .O(N__18919),
            .I(N__18915));
    SRMux I__3583 (
            .O(N__18918),
            .I(N__18912));
    LocalMux I__3582 (
            .O(N__18915),
            .I(N__18909));
    LocalMux I__3581 (
            .O(N__18912),
            .I(N__18906));
    Span4Mux_h I__3580 (
            .O(N__18909),
            .I(N__18903));
    Odrv12 I__3579 (
            .O(N__18906),
            .I(\uu2.vram_wr_en_0_iZ0 ));
    Odrv4 I__3578 (
            .O(N__18903),
            .I(\uu2.vram_wr_en_0_iZ0 ));
    InMux I__3577 (
            .O(N__18898),
            .I(N__18895));
    LocalMux I__3576 (
            .O(N__18895),
            .I(\uu2.un1_w_user_lf_0 ));
    CascadeMux I__3575 (
            .O(N__18892),
            .I(N__18888));
    InMux I__3574 (
            .O(N__18891),
            .I(N__18883));
    InMux I__3573 (
            .O(N__18888),
            .I(N__18883));
    LocalMux I__3572 (
            .O(N__18883),
            .I(\uu2.un3_w_addr_user ));
    InMux I__3571 (
            .O(N__18880),
            .I(N__18871));
    InMux I__3570 (
            .O(N__18879),
            .I(N__18871));
    InMux I__3569 (
            .O(N__18878),
            .I(N__18871));
    LocalMux I__3568 (
            .O(N__18871),
            .I(\uu2.un1_w_user_cr_0 ));
    CascadeMux I__3567 (
            .O(N__18868),
            .I(\uu2.un1_w_user_cr_0_cascade_ ));
    InMux I__3566 (
            .O(N__18865),
            .I(N__18858));
    InMux I__3565 (
            .O(N__18864),
            .I(N__18858));
    InMux I__3564 (
            .O(N__18863),
            .I(N__18855));
    LocalMux I__3563 (
            .O(N__18858),
            .I(N__18852));
    LocalMux I__3562 (
            .O(N__18855),
            .I(\uu2.N_71 ));
    Odrv12 I__3561 (
            .O(N__18852),
            .I(\uu2.N_71 ));
    CascadeMux I__3560 (
            .O(N__18847),
            .I(\uu2.un4_w_user_data_rdyZ0Z_0_cascade_ ));
    InMux I__3559 (
            .O(N__18844),
            .I(N__18841));
    LocalMux I__3558 (
            .O(N__18841),
            .I(N__18838));
    Span4Mux_s3_h I__3557 (
            .O(N__18838),
            .I(N__18835));
    Span4Mux_h I__3556 (
            .O(N__18835),
            .I(N__18832));
    Odrv4 I__3555 (
            .O(N__18832),
            .I(\uu2.mem0.w_data_6 ));
    InMux I__3554 (
            .O(N__18829),
            .I(N__18826));
    LocalMux I__3553 (
            .O(N__18826),
            .I(\uu2.un1_w_user_crZ0Z_4 ));
    InMux I__3552 (
            .O(N__18823),
            .I(N__18820));
    LocalMux I__3551 (
            .O(N__18820),
            .I(\uu2.un1_w_user_lfZ0Z_4 ));
    InMux I__3550 (
            .O(N__18817),
            .I(N__18814));
    LocalMux I__3549 (
            .O(N__18814),
            .I(N__18811));
    Span4Mux_s3_h I__3548 (
            .O(N__18811),
            .I(N__18808));
    Span4Mux_h I__3547 (
            .O(N__18808),
            .I(N__18805));
    Odrv4 I__3546 (
            .O(N__18805),
            .I(\uu2.mem0.w_data_2 ));
    InMux I__3545 (
            .O(N__18802),
            .I(N__18787));
    InMux I__3544 (
            .O(N__18801),
            .I(N__18787));
    InMux I__3543 (
            .O(N__18800),
            .I(N__18787));
    InMux I__3542 (
            .O(N__18799),
            .I(N__18787));
    InMux I__3541 (
            .O(N__18798),
            .I(N__18787));
    LocalMux I__3540 (
            .O(N__18787),
            .I(N__18782));
    InMux I__3539 (
            .O(N__18786),
            .I(N__18779));
    InMux I__3538 (
            .O(N__18785),
            .I(N__18776));
    Span4Mux_v I__3537 (
            .O(N__18782),
            .I(N__18764));
    LocalMux I__3536 (
            .O(N__18779),
            .I(N__18764));
    LocalMux I__3535 (
            .O(N__18776),
            .I(N__18764));
    InMux I__3534 (
            .O(N__18775),
            .I(N__18761));
    InMux I__3533 (
            .O(N__18774),
            .I(N__18752));
    InMux I__3532 (
            .O(N__18773),
            .I(N__18752));
    InMux I__3531 (
            .O(N__18772),
            .I(N__18752));
    InMux I__3530 (
            .O(N__18771),
            .I(N__18752));
    Span4Mux_h I__3529 (
            .O(N__18764),
            .I(N__18745));
    LocalMux I__3528 (
            .O(N__18761),
            .I(N__18742));
    LocalMux I__3527 (
            .O(N__18752),
            .I(N__18739));
    InMux I__3526 (
            .O(N__18751),
            .I(N__18734));
    InMux I__3525 (
            .O(N__18750),
            .I(N__18734));
    InMux I__3524 (
            .O(N__18749),
            .I(N__18731));
    InMux I__3523 (
            .O(N__18748),
            .I(N__18728));
    Odrv4 I__3522 (
            .O(N__18745),
            .I(\uu2.un4_w_user_data_rdyZ0Z_0 ));
    Odrv12 I__3521 (
            .O(N__18742),
            .I(\uu2.un4_w_user_data_rdyZ0Z_0 ));
    Odrv4 I__3520 (
            .O(N__18739),
            .I(\uu2.un4_w_user_data_rdyZ0Z_0 ));
    LocalMux I__3519 (
            .O(N__18734),
            .I(\uu2.un4_w_user_data_rdyZ0Z_0 ));
    LocalMux I__3518 (
            .O(N__18731),
            .I(\uu2.un4_w_user_data_rdyZ0Z_0 ));
    LocalMux I__3517 (
            .O(N__18728),
            .I(\uu2.un4_w_user_data_rdyZ0Z_0 ));
    CascadeMux I__3516 (
            .O(N__18715),
            .I(N__18712));
    InMux I__3515 (
            .O(N__18712),
            .I(N__18709));
    LocalMux I__3514 (
            .O(N__18709),
            .I(N__18706));
    Span12Mux_s7_h I__3513 (
            .O(N__18706),
            .I(N__18703));
    Odrv12 I__3512 (
            .O(N__18703),
            .I(\uu2.mem0.w_addr_0 ));
    CascadeMux I__3511 (
            .O(N__18700),
            .I(\Lab_UT.uu0.un4_l_count_14_cascade_ ));
    CascadeMux I__3510 (
            .O(N__18697),
            .I(\Lab_UT.uu0.un187_ci_1_cascade_ ));
    CascadeMux I__3509 (
            .O(N__18694),
            .I(N__18691));
    InMux I__3508 (
            .O(N__18691),
            .I(N__18685));
    InMux I__3507 (
            .O(N__18690),
            .I(N__18678));
    InMux I__3506 (
            .O(N__18689),
            .I(N__18678));
    InMux I__3505 (
            .O(N__18688),
            .I(N__18678));
    LocalMux I__3504 (
            .O(N__18685),
            .I(\Lab_UT.uu0.un154_ci_9 ));
    LocalMux I__3503 (
            .O(N__18678),
            .I(\Lab_UT.uu0.un154_ci_9 ));
    CascadeMux I__3502 (
            .O(N__18673),
            .I(N__18667));
    CascadeMux I__3501 (
            .O(N__18672),
            .I(N__18664));
    CascadeMux I__3500 (
            .O(N__18671),
            .I(N__18661));
    InMux I__3499 (
            .O(N__18670),
            .I(N__18656));
    InMux I__3498 (
            .O(N__18667),
            .I(N__18656));
    InMux I__3497 (
            .O(N__18664),
            .I(N__18651));
    InMux I__3496 (
            .O(N__18661),
            .I(N__18651));
    LocalMux I__3495 (
            .O(N__18656),
            .I(\Lab_UT.uu0.l_countZ0Z_14 ));
    LocalMux I__3494 (
            .O(N__18651),
            .I(\Lab_UT.uu0.l_countZ0Z_14 ));
    InMux I__3493 (
            .O(N__18646),
            .I(N__18640));
    InMux I__3492 (
            .O(N__18645),
            .I(N__18633));
    InMux I__3491 (
            .O(N__18644),
            .I(N__18633));
    InMux I__3490 (
            .O(N__18643),
            .I(N__18633));
    LocalMux I__3489 (
            .O(N__18640),
            .I(N__18628));
    LocalMux I__3488 (
            .O(N__18633),
            .I(N__18628));
    Span4Mux_h I__3487 (
            .O(N__18628),
            .I(N__18625));
    Odrv4 I__3486 (
            .O(N__18625),
            .I(\Lab_UT.uu0.un4_l_count_0_8 ));
    InMux I__3485 (
            .O(N__18622),
            .I(N__18613));
    InMux I__3484 (
            .O(N__18621),
            .I(N__18613));
    InMux I__3483 (
            .O(N__18620),
            .I(N__18613));
    LocalMux I__3482 (
            .O(N__18613),
            .I(\Lab_UT.uu0.un198_ci_2 ));
    CascadeMux I__3481 (
            .O(N__18610),
            .I(N__18605));
    CascadeMux I__3480 (
            .O(N__18609),
            .I(N__18598));
    CascadeMux I__3479 (
            .O(N__18608),
            .I(N__18595));
    InMux I__3478 (
            .O(N__18605),
            .I(N__18585));
    InMux I__3477 (
            .O(N__18604),
            .I(N__18585));
    InMux I__3476 (
            .O(N__18603),
            .I(N__18585));
    InMux I__3475 (
            .O(N__18602),
            .I(N__18582));
    InMux I__3474 (
            .O(N__18601),
            .I(N__18577));
    InMux I__3473 (
            .O(N__18598),
            .I(N__18577));
    InMux I__3472 (
            .O(N__18595),
            .I(N__18568));
    InMux I__3471 (
            .O(N__18594),
            .I(N__18568));
    InMux I__3470 (
            .O(N__18593),
            .I(N__18568));
    InMux I__3469 (
            .O(N__18592),
            .I(N__18568));
    LocalMux I__3468 (
            .O(N__18585),
            .I(\Lab_UT.uu0.un110_ci ));
    LocalMux I__3467 (
            .O(N__18582),
            .I(\Lab_UT.uu0.un110_ci ));
    LocalMux I__3466 (
            .O(N__18577),
            .I(\Lab_UT.uu0.un110_ci ));
    LocalMux I__3465 (
            .O(N__18568),
            .I(\Lab_UT.uu0.un110_ci ));
    InMux I__3464 (
            .O(N__18559),
            .I(N__18547));
    InMux I__3463 (
            .O(N__18558),
            .I(N__18547));
    InMux I__3462 (
            .O(N__18557),
            .I(N__18547));
    InMux I__3461 (
            .O(N__18556),
            .I(N__18540));
    InMux I__3460 (
            .O(N__18555),
            .I(N__18540));
    InMux I__3459 (
            .O(N__18554),
            .I(N__18540));
    LocalMux I__3458 (
            .O(N__18547),
            .I(\Lab_UT.uu0.l_countZ0Z_8 ));
    LocalMux I__3457 (
            .O(N__18540),
            .I(\Lab_UT.uu0.l_countZ0Z_8 ));
    CEMux I__3456 (
            .O(N__18535),
            .I(N__18532));
    LocalMux I__3455 (
            .O(N__18532),
            .I(N__18529));
    Span4Mux_s2_v I__3454 (
            .O(N__18529),
            .I(N__18526));
    Odrv4 I__3453 (
            .O(N__18526),
            .I(\uu2.un28_w_addr_user_i_0 ));
    CascadeMux I__3452 (
            .O(N__18523),
            .I(\uu2.un1_w_user_lf_0_cascade_ ));
    CascadeMux I__3451 (
            .O(N__18520),
            .I(\Lab_UT.uu0.un99_ci_0_cascade_ ));
    CascadeMux I__3450 (
            .O(N__18517),
            .I(N__18514));
    InMux I__3449 (
            .O(N__18514),
            .I(N__18508));
    InMux I__3448 (
            .O(N__18513),
            .I(N__18508));
    LocalMux I__3447 (
            .O(N__18508),
            .I(\Lab_UT.uu0.un88_ci_3 ));
    CascadeMux I__3446 (
            .O(N__18505),
            .I(\Lab_UT.uu0.un88_ci_3_cascade_ ));
    InMux I__3445 (
            .O(N__18502),
            .I(N__18495));
    InMux I__3444 (
            .O(N__18501),
            .I(N__18495));
    InMux I__3443 (
            .O(N__18500),
            .I(N__18492));
    LocalMux I__3442 (
            .O(N__18495),
            .I(\Lab_UT.uu0.l_countZ0Z_7 ));
    LocalMux I__3441 (
            .O(N__18492),
            .I(\Lab_UT.uu0.l_countZ0Z_7 ));
    CascadeMux I__3440 (
            .O(N__18487),
            .I(N__18483));
    CascadeMux I__3439 (
            .O(N__18486),
            .I(N__18480));
    InMux I__3438 (
            .O(N__18483),
            .I(N__18476));
    InMux I__3437 (
            .O(N__18480),
            .I(N__18471));
    InMux I__3436 (
            .O(N__18479),
            .I(N__18471));
    LocalMux I__3435 (
            .O(N__18476),
            .I(N__18468));
    LocalMux I__3434 (
            .O(N__18471),
            .I(\Lab_UT.uu0.l_countZ0Z_17 ));
    Odrv4 I__3433 (
            .O(N__18468),
            .I(\Lab_UT.uu0.l_countZ0Z_17 ));
    CascadeMux I__3432 (
            .O(N__18463),
            .I(\Lab_UT.uu0.un110_ci_cascade_ ));
    InMux I__3431 (
            .O(N__18460),
            .I(N__18457));
    LocalMux I__3430 (
            .O(N__18457),
            .I(\Lab_UT.uu0.un220_ci ));
    InMux I__3429 (
            .O(N__18454),
            .I(N__18447));
    InMux I__3428 (
            .O(N__18453),
            .I(N__18440));
    InMux I__3427 (
            .O(N__18452),
            .I(N__18440));
    InMux I__3426 (
            .O(N__18451),
            .I(N__18440));
    InMux I__3425 (
            .O(N__18450),
            .I(N__18437));
    LocalMux I__3424 (
            .O(N__18447),
            .I(\Lab_UT.uu0.l_countZ0Z_9 ));
    LocalMux I__3423 (
            .O(N__18440),
            .I(\Lab_UT.uu0.l_countZ0Z_9 ));
    LocalMux I__3422 (
            .O(N__18437),
            .I(\Lab_UT.uu0.l_countZ0Z_9 ));
    InMux I__3421 (
            .O(N__18430),
            .I(N__18424));
    InMux I__3420 (
            .O(N__18429),
            .I(N__18421));
    InMux I__3419 (
            .O(N__18428),
            .I(N__18416));
    InMux I__3418 (
            .O(N__18427),
            .I(N__18416));
    LocalMux I__3417 (
            .O(N__18424),
            .I(\Lab_UT.uu0.l_countZ0Z_10 ));
    LocalMux I__3416 (
            .O(N__18421),
            .I(\Lab_UT.uu0.l_countZ0Z_10 ));
    LocalMux I__3415 (
            .O(N__18416),
            .I(\Lab_UT.uu0.l_countZ0Z_10 ));
    InMux I__3414 (
            .O(N__18409),
            .I(N__18406));
    LocalMux I__3413 (
            .O(N__18406),
            .I(N__18403));
    Odrv4 I__3412 (
            .O(N__18403),
            .I(\Lab_UT.dictrl.decoder.g0_3Z0Z_0 ));
    CascadeMux I__3411 (
            .O(N__18400),
            .I(N__18397));
    InMux I__3410 (
            .O(N__18397),
            .I(N__18394));
    LocalMux I__3409 (
            .O(N__18394),
            .I(N__18391));
    Span4Mux_h I__3408 (
            .O(N__18391),
            .I(N__18388));
    Odrv4 I__3407 (
            .O(N__18388),
            .I(\Lab_UT.dictrl.de_cr_1_2 ));
    InMux I__3406 (
            .O(N__18385),
            .I(N__18382));
    LocalMux I__3405 (
            .O(N__18382),
            .I(\Lab_UT.dictrl.decoder.g0_4Z0Z_3 ));
    CascadeMux I__3404 (
            .O(N__18379),
            .I(\Lab_UT.dictrl.decoder.g0_3_2_cascade_ ));
    CascadeMux I__3403 (
            .O(N__18376),
            .I(N__18372));
    InMux I__3402 (
            .O(N__18375),
            .I(N__18368));
    InMux I__3401 (
            .O(N__18372),
            .I(N__18361));
    InMux I__3400 (
            .O(N__18371),
            .I(N__18361));
    LocalMux I__3399 (
            .O(N__18368),
            .I(N__18358));
    InMux I__3398 (
            .O(N__18367),
            .I(N__18353));
    InMux I__3397 (
            .O(N__18366),
            .I(N__18353));
    LocalMux I__3396 (
            .O(N__18361),
            .I(N__18348));
    Span4Mux_h I__3395 (
            .O(N__18358),
            .I(N__18348));
    LocalMux I__3394 (
            .O(N__18353),
            .I(Lab_UT_dictrl_decoder_de_cr_1_1));
    Odrv4 I__3393 (
            .O(N__18348),
            .I(Lab_UT_dictrl_decoder_de_cr_1_1));
    CascadeMux I__3392 (
            .O(N__18343),
            .I(N__18340));
    InMux I__3391 (
            .O(N__18340),
            .I(N__18337));
    LocalMux I__3390 (
            .O(N__18337),
            .I(N__18334));
    Odrv4 I__3389 (
            .O(N__18334),
            .I(\Lab_UT.dictrl.de_cr_2_0 ));
    CascadeMux I__3388 (
            .O(N__18331),
            .I(N__18328));
    InMux I__3387 (
            .O(N__18328),
            .I(N__18325));
    LocalMux I__3386 (
            .O(N__18325),
            .I(\Lab_UT.dictrl.decoder.g0_4_1 ));
    CascadeMux I__3385 (
            .O(N__18322),
            .I(N__18314));
    CascadeMux I__3384 (
            .O(N__18321),
            .I(N__18311));
    CascadeMux I__3383 (
            .O(N__18320),
            .I(N__18308));
    InMux I__3382 (
            .O(N__18319),
            .I(N__18301));
    InMux I__3381 (
            .O(N__18318),
            .I(N__18301));
    InMux I__3380 (
            .O(N__18317),
            .I(N__18294));
    InMux I__3379 (
            .O(N__18314),
            .I(N__18294));
    InMux I__3378 (
            .O(N__18311),
            .I(N__18294));
    InMux I__3377 (
            .O(N__18308),
            .I(N__18287));
    InMux I__3376 (
            .O(N__18307),
            .I(N__18287));
    InMux I__3375 (
            .O(N__18306),
            .I(N__18287));
    LocalMux I__3374 (
            .O(N__18301),
            .I(buart__rx_bitcount_4));
    LocalMux I__3373 (
            .O(N__18294),
            .I(buart__rx_bitcount_4));
    LocalMux I__3372 (
            .O(N__18287),
            .I(buart__rx_bitcount_4));
    InMux I__3371 (
            .O(N__18280),
            .I(N__18275));
    InMux I__3370 (
            .O(N__18279),
            .I(N__18264));
    InMux I__3369 (
            .O(N__18278),
            .I(N__18264));
    LocalMux I__3368 (
            .O(N__18275),
            .I(N__18261));
    InMux I__3367 (
            .O(N__18274),
            .I(N__18254));
    InMux I__3366 (
            .O(N__18273),
            .I(N__18254));
    InMux I__3365 (
            .O(N__18272),
            .I(N__18254));
    InMux I__3364 (
            .O(N__18271),
            .I(N__18247));
    InMux I__3363 (
            .O(N__18270),
            .I(N__18247));
    InMux I__3362 (
            .O(N__18269),
            .I(N__18247));
    LocalMux I__3361 (
            .O(N__18264),
            .I(buart__rx_bitcount_3));
    Odrv4 I__3360 (
            .O(N__18261),
            .I(buart__rx_bitcount_3));
    LocalMux I__3359 (
            .O(N__18254),
            .I(buart__rx_bitcount_3));
    LocalMux I__3358 (
            .O(N__18247),
            .I(buart__rx_bitcount_3));
    InMux I__3357 (
            .O(N__18238),
            .I(N__18227));
    InMux I__3356 (
            .O(N__18237),
            .I(N__18227));
    InMux I__3355 (
            .O(N__18236),
            .I(N__18217));
    InMux I__3354 (
            .O(N__18235),
            .I(N__18217));
    InMux I__3353 (
            .O(N__18234),
            .I(N__18217));
    InMux I__3352 (
            .O(N__18233),
            .I(N__18212));
    InMux I__3351 (
            .O(N__18232),
            .I(N__18212));
    LocalMux I__3350 (
            .O(N__18227),
            .I(N__18209));
    InMux I__3349 (
            .O(N__18226),
            .I(N__18204));
    InMux I__3348 (
            .O(N__18225),
            .I(N__18204));
    InMux I__3347 (
            .O(N__18224),
            .I(N__18201));
    LocalMux I__3346 (
            .O(N__18217),
            .I(buart__rx_bitcount_2));
    LocalMux I__3345 (
            .O(N__18212),
            .I(buart__rx_bitcount_2));
    Odrv4 I__3344 (
            .O(N__18209),
            .I(buart__rx_bitcount_2));
    LocalMux I__3343 (
            .O(N__18204),
            .I(buart__rx_bitcount_2));
    LocalMux I__3342 (
            .O(N__18201),
            .I(buart__rx_bitcount_2));
    CascadeMux I__3341 (
            .O(N__18190),
            .I(\Lab_UT.dictrl.g0_8_cascade_ ));
    InMux I__3340 (
            .O(N__18187),
            .I(N__18183));
    CascadeMux I__3339 (
            .O(N__18186),
            .I(N__18180));
    LocalMux I__3338 (
            .O(N__18183),
            .I(N__18176));
    InMux I__3337 (
            .O(N__18180),
            .I(N__18168));
    InMux I__3336 (
            .O(N__18179),
            .I(N__18165));
    Span4Mux_v I__3335 (
            .O(N__18176),
            .I(N__18162));
    InMux I__3334 (
            .O(N__18175),
            .I(N__18155));
    InMux I__3333 (
            .O(N__18174),
            .I(N__18155));
    InMux I__3332 (
            .O(N__18173),
            .I(N__18155));
    InMux I__3331 (
            .O(N__18172),
            .I(N__18152));
    InMux I__3330 (
            .O(N__18171),
            .I(N__18149));
    LocalMux I__3329 (
            .O(N__18168),
            .I(N__18146));
    LocalMux I__3328 (
            .O(N__18165),
            .I(N__18143));
    Odrv4 I__3327 (
            .O(N__18162),
            .I(buart__rx_valid_2_0));
    LocalMux I__3326 (
            .O(N__18155),
            .I(buart__rx_valid_2_0));
    LocalMux I__3325 (
            .O(N__18152),
            .I(buart__rx_valid_2_0));
    LocalMux I__3324 (
            .O(N__18149),
            .I(buart__rx_valid_2_0));
    Odrv4 I__3323 (
            .O(N__18146),
            .I(buart__rx_valid_2_0));
    Odrv4 I__3322 (
            .O(N__18143),
            .I(buart__rx_valid_2_0));
    InMux I__3321 (
            .O(N__18130),
            .I(N__18127));
    LocalMux I__3320 (
            .O(N__18127),
            .I(N__18124));
    Span4Mux_h I__3319 (
            .O(N__18124),
            .I(N__18121));
    Span4Mux_v I__3318 (
            .O(N__18121),
            .I(N__18118));
    Odrv4 I__3317 (
            .O(N__18118),
            .I(\Lab_UT.dictrl.g0_11 ));
    InMux I__3316 (
            .O(N__18115),
            .I(N__18112));
    LocalMux I__3315 (
            .O(N__18112),
            .I(N__18108));
    InMux I__3314 (
            .O(N__18111),
            .I(N__18105));
    Span4Mux_v I__3313 (
            .O(N__18108),
            .I(N__18102));
    LocalMux I__3312 (
            .O(N__18105),
            .I(N__18099));
    Span4Mux_h I__3311 (
            .O(N__18102),
            .I(N__18096));
    Span4Mux_h I__3310 (
            .O(N__18099),
            .I(N__18093));
    Odrv4 I__3309 (
            .O(N__18096),
            .I(\Lab_UT.dictrl.currState_2_RNIEPCJZ0Z_1 ));
    Odrv4 I__3308 (
            .O(N__18093),
            .I(\Lab_UT.dictrl.currState_2_RNIEPCJZ0Z_1 ));
    InMux I__3307 (
            .O(N__18088),
            .I(N__18085));
    LocalMux I__3306 (
            .O(N__18085),
            .I(N__18081));
    InMux I__3305 (
            .O(N__18084),
            .I(N__18078));
    Span4Mux_h I__3304 (
            .O(N__18081),
            .I(N__18075));
    LocalMux I__3303 (
            .O(N__18078),
            .I(\Lab_UT.dictrl.nextState_0_3 ));
    Odrv4 I__3302 (
            .O(N__18075),
            .I(\Lab_UT.dictrl.nextState_0_3 ));
    InMux I__3301 (
            .O(N__18070),
            .I(N__18067));
    LocalMux I__3300 (
            .O(N__18067),
            .I(\Lab_UT.dictrl.N_1612_0 ));
    InMux I__3299 (
            .O(N__18064),
            .I(N__18048));
    InMux I__3298 (
            .O(N__18063),
            .I(N__18048));
    InMux I__3297 (
            .O(N__18062),
            .I(N__18043));
    InMux I__3296 (
            .O(N__18061),
            .I(N__18038));
    InMux I__3295 (
            .O(N__18060),
            .I(N__18031));
    InMux I__3294 (
            .O(N__18059),
            .I(N__18031));
    InMux I__3293 (
            .O(N__18058),
            .I(N__18031));
    InMux I__3292 (
            .O(N__18057),
            .I(N__18026));
    InMux I__3291 (
            .O(N__18056),
            .I(N__18026));
    InMux I__3290 (
            .O(N__18055),
            .I(N__18023));
    InMux I__3289 (
            .O(N__18054),
            .I(N__18018));
    InMux I__3288 (
            .O(N__18053),
            .I(N__18018));
    LocalMux I__3287 (
            .O(N__18048),
            .I(N__18015));
    CascadeMux I__3286 (
            .O(N__18047),
            .I(N__18010));
    InMux I__3285 (
            .O(N__18046),
            .I(N__18003));
    LocalMux I__3284 (
            .O(N__18043),
            .I(N__18000));
    InMux I__3283 (
            .O(N__18042),
            .I(N__17997));
    InMux I__3282 (
            .O(N__18041),
            .I(N__17994));
    LocalMux I__3281 (
            .O(N__18038),
            .I(N__17987));
    LocalMux I__3280 (
            .O(N__18031),
            .I(N__17987));
    LocalMux I__3279 (
            .O(N__18026),
            .I(N__17987));
    LocalMux I__3278 (
            .O(N__18023),
            .I(N__17982));
    LocalMux I__3277 (
            .O(N__18018),
            .I(N__17982));
    Span4Mux_v I__3276 (
            .O(N__18015),
            .I(N__17979));
    InMux I__3275 (
            .O(N__18014),
            .I(N__17976));
    InMux I__3274 (
            .O(N__18013),
            .I(N__17973));
    InMux I__3273 (
            .O(N__18010),
            .I(N__17966));
    InMux I__3272 (
            .O(N__18009),
            .I(N__17966));
    InMux I__3271 (
            .O(N__18008),
            .I(N__17966));
    InMux I__3270 (
            .O(N__18007),
            .I(N__17963));
    InMux I__3269 (
            .O(N__18006),
            .I(N__17960));
    LocalMux I__3268 (
            .O(N__18003),
            .I(N__17951));
    Span4Mux_h I__3267 (
            .O(N__18000),
            .I(N__17951));
    LocalMux I__3266 (
            .O(N__17997),
            .I(N__17951));
    LocalMux I__3265 (
            .O(N__17994),
            .I(N__17951));
    Span4Mux_v I__3264 (
            .O(N__17987),
            .I(N__17946));
    Span4Mux_v I__3263 (
            .O(N__17982),
            .I(N__17946));
    Odrv4 I__3262 (
            .O(N__17979),
            .I(\Lab_UT.dictrl.currState_2_RNI2P2AZ0Z_2 ));
    LocalMux I__3261 (
            .O(N__17976),
            .I(\Lab_UT.dictrl.currState_2_RNI2P2AZ0Z_2 ));
    LocalMux I__3260 (
            .O(N__17973),
            .I(\Lab_UT.dictrl.currState_2_RNI2P2AZ0Z_2 ));
    LocalMux I__3259 (
            .O(N__17966),
            .I(\Lab_UT.dictrl.currState_2_RNI2P2AZ0Z_2 ));
    LocalMux I__3258 (
            .O(N__17963),
            .I(\Lab_UT.dictrl.currState_2_RNI2P2AZ0Z_2 ));
    LocalMux I__3257 (
            .O(N__17960),
            .I(\Lab_UT.dictrl.currState_2_RNI2P2AZ0Z_2 ));
    Odrv4 I__3256 (
            .O(N__17951),
            .I(\Lab_UT.dictrl.currState_2_RNI2P2AZ0Z_2 ));
    Odrv4 I__3255 (
            .O(N__17946),
            .I(\Lab_UT.dictrl.currState_2_RNI2P2AZ0Z_2 ));
    CascadeMux I__3254 (
            .O(N__17929),
            .I(N__17921));
    InMux I__3253 (
            .O(N__17928),
            .I(N__17907));
    InMux I__3252 (
            .O(N__17927),
            .I(N__17895));
    InMux I__3251 (
            .O(N__17926),
            .I(N__17895));
    InMux I__3250 (
            .O(N__17925),
            .I(N__17895));
    InMux I__3249 (
            .O(N__17924),
            .I(N__17895));
    InMux I__3248 (
            .O(N__17921),
            .I(N__17889));
    InMux I__3247 (
            .O(N__17920),
            .I(N__17883));
    InMux I__3246 (
            .O(N__17919),
            .I(N__17876));
    InMux I__3245 (
            .O(N__17918),
            .I(N__17876));
    InMux I__3244 (
            .O(N__17917),
            .I(N__17876));
    InMux I__3243 (
            .O(N__17916),
            .I(N__17873));
    InMux I__3242 (
            .O(N__17915),
            .I(N__17870));
    InMux I__3241 (
            .O(N__17914),
            .I(N__17863));
    InMux I__3240 (
            .O(N__17913),
            .I(N__17863));
    InMux I__3239 (
            .O(N__17912),
            .I(N__17863));
    InMux I__3238 (
            .O(N__17911),
            .I(N__17856));
    CascadeMux I__3237 (
            .O(N__17910),
            .I(N__17851));
    LocalMux I__3236 (
            .O(N__17907),
            .I(N__17848));
    InMux I__3235 (
            .O(N__17906),
            .I(N__17841));
    InMux I__3234 (
            .O(N__17905),
            .I(N__17841));
    InMux I__3233 (
            .O(N__17904),
            .I(N__17841));
    LocalMux I__3232 (
            .O(N__17895),
            .I(N__17838));
    CascadeMux I__3231 (
            .O(N__17894),
            .I(N__17835));
    CascadeMux I__3230 (
            .O(N__17893),
            .I(N__17832));
    CascadeMux I__3229 (
            .O(N__17892),
            .I(N__17829));
    LocalMux I__3228 (
            .O(N__17889),
            .I(N__17825));
    InMux I__3227 (
            .O(N__17888),
            .I(N__17818));
    InMux I__3226 (
            .O(N__17887),
            .I(N__17818));
    InMux I__3225 (
            .O(N__17886),
            .I(N__17818));
    LocalMux I__3224 (
            .O(N__17883),
            .I(N__17811));
    LocalMux I__3223 (
            .O(N__17876),
            .I(N__17811));
    LocalMux I__3222 (
            .O(N__17873),
            .I(N__17811));
    LocalMux I__3221 (
            .O(N__17870),
            .I(N__17806));
    LocalMux I__3220 (
            .O(N__17863),
            .I(N__17806));
    InMux I__3219 (
            .O(N__17862),
            .I(N__17803));
    InMux I__3218 (
            .O(N__17861),
            .I(N__17800));
    InMux I__3217 (
            .O(N__17860),
            .I(N__17795));
    InMux I__3216 (
            .O(N__17859),
            .I(N__17795));
    LocalMux I__3215 (
            .O(N__17856),
            .I(N__17792));
    InMux I__3214 (
            .O(N__17855),
            .I(N__17785));
    InMux I__3213 (
            .O(N__17854),
            .I(N__17785));
    InMux I__3212 (
            .O(N__17851),
            .I(N__17785));
    Span4Mux_v I__3211 (
            .O(N__17848),
            .I(N__17778));
    LocalMux I__3210 (
            .O(N__17841),
            .I(N__17778));
    Span4Mux_v I__3209 (
            .O(N__17838),
            .I(N__17778));
    InMux I__3208 (
            .O(N__17835),
            .I(N__17773));
    InMux I__3207 (
            .O(N__17832),
            .I(N__17773));
    InMux I__3206 (
            .O(N__17829),
            .I(N__17770));
    InMux I__3205 (
            .O(N__17828),
            .I(N__17767));
    Span4Mux_v I__3204 (
            .O(N__17825),
            .I(N__17760));
    LocalMux I__3203 (
            .O(N__17818),
            .I(N__17760));
    Span4Mux_v I__3202 (
            .O(N__17811),
            .I(N__17760));
    Span4Mux_h I__3201 (
            .O(N__17806),
            .I(N__17753));
    LocalMux I__3200 (
            .O(N__17803),
            .I(N__17753));
    LocalMux I__3199 (
            .O(N__17800),
            .I(N__17753));
    LocalMux I__3198 (
            .O(N__17795),
            .I(N__17750));
    Span12Mux_s10_h I__3197 (
            .O(N__17792),
            .I(N__17745));
    LocalMux I__3196 (
            .O(N__17785),
            .I(N__17745));
    Span4Mux_h I__3195 (
            .O(N__17778),
            .I(N__17742));
    LocalMux I__3194 (
            .O(N__17773),
            .I(Lab_UT_dictrl_currState_1));
    LocalMux I__3193 (
            .O(N__17770),
            .I(Lab_UT_dictrl_currState_1));
    LocalMux I__3192 (
            .O(N__17767),
            .I(Lab_UT_dictrl_currState_1));
    Odrv4 I__3191 (
            .O(N__17760),
            .I(Lab_UT_dictrl_currState_1));
    Odrv4 I__3190 (
            .O(N__17753),
            .I(Lab_UT_dictrl_currState_1));
    Odrv4 I__3189 (
            .O(N__17750),
            .I(Lab_UT_dictrl_currState_1));
    Odrv12 I__3188 (
            .O(N__17745),
            .I(Lab_UT_dictrl_currState_1));
    Odrv4 I__3187 (
            .O(N__17742),
            .I(Lab_UT_dictrl_currState_1));
    InMux I__3186 (
            .O(N__17725),
            .I(N__17721));
    InMux I__3185 (
            .O(N__17724),
            .I(N__17718));
    LocalMux I__3184 (
            .O(N__17721),
            .I(N__17713));
    LocalMux I__3183 (
            .O(N__17718),
            .I(N__17713));
    Odrv12 I__3182 (
            .O(N__17713),
            .I(\Lab_UT.dictrl.G_19_0_a7_2 ));
    InMux I__3181 (
            .O(N__17710),
            .I(N__17707));
    LocalMux I__3180 (
            .O(N__17707),
            .I(N__17704));
    Odrv4 I__3179 (
            .O(N__17704),
            .I(\Lab_UT.dictrl.decoder.g0_2Z0Z_2 ));
    CascadeMux I__3178 (
            .O(N__17701),
            .I(Lab_UT_dictrl_decoder_de_cr_2_cascade_));
    InMux I__3177 (
            .O(N__17698),
            .I(N__17691));
    InMux I__3176 (
            .O(N__17697),
            .I(N__17688));
    InMux I__3175 (
            .O(N__17696),
            .I(N__17683));
    InMux I__3174 (
            .O(N__17695),
            .I(N__17683));
    InMux I__3173 (
            .O(N__17694),
            .I(N__17680));
    LocalMux I__3172 (
            .O(N__17691),
            .I(buart__rx_bitcount_2_rep1));
    LocalMux I__3171 (
            .O(N__17688),
            .I(buart__rx_bitcount_2_rep1));
    LocalMux I__3170 (
            .O(N__17683),
            .I(buart__rx_bitcount_2_rep1));
    LocalMux I__3169 (
            .O(N__17680),
            .I(buart__rx_bitcount_2_rep1));
    CascadeMux I__3168 (
            .O(N__17671),
            .I(\Lab_UT.dictrl.decoder.g0_4_0_cascade_ ));
    InMux I__3167 (
            .O(N__17668),
            .I(N__17664));
    InMux I__3166 (
            .O(N__17667),
            .I(N__17661));
    LocalMux I__3165 (
            .O(N__17664),
            .I(N__17657));
    LocalMux I__3164 (
            .O(N__17661),
            .I(N__17654));
    InMux I__3163 (
            .O(N__17660),
            .I(N__17651));
    Span4Mux_s3_h I__3162 (
            .O(N__17657),
            .I(N__17642));
    Span4Mux_s3_v I__3161 (
            .O(N__17654),
            .I(N__17642));
    LocalMux I__3160 (
            .O(N__17651),
            .I(N__17642));
    InMux I__3159 (
            .O(N__17650),
            .I(N__17639));
    InMux I__3158 (
            .O(N__17649),
            .I(N__17636));
    Odrv4 I__3157 (
            .O(N__17642),
            .I(\Lab_UT.dictrl.de_cr_1_0 ));
    LocalMux I__3156 (
            .O(N__17639),
            .I(\Lab_UT.dictrl.de_cr_1_0 ));
    LocalMux I__3155 (
            .O(N__17636),
            .I(\Lab_UT.dictrl.de_cr_1_0 ));
    InMux I__3154 (
            .O(N__17629),
            .I(N__17626));
    LocalMux I__3153 (
            .O(N__17626),
            .I(N__17623));
    Span4Mux_h I__3152 (
            .O(N__17623),
            .I(N__17620));
    Odrv4 I__3151 (
            .O(N__17620),
            .I(\Lab_UT.dictrl.de_cr_0 ));
    InMux I__3150 (
            .O(N__17617),
            .I(N__17613));
    InMux I__3149 (
            .O(N__17616),
            .I(N__17610));
    LocalMux I__3148 (
            .O(N__17613),
            .I(N__17607));
    LocalMux I__3147 (
            .O(N__17610),
            .I(bu_rx_data_fast_2));
    Odrv4 I__3146 (
            .O(N__17607),
            .I(bu_rx_data_fast_2));
    CascadeMux I__3145 (
            .O(N__17602),
            .I(\Lab_UT.dictrl.r_dicLdMtens15_1i_cascade_ ));
    InMux I__3144 (
            .O(N__17599),
            .I(N__17596));
    LocalMux I__3143 (
            .O(N__17596),
            .I(N__17593));
    Span4Mux_h I__3142 (
            .O(N__17593),
            .I(N__17590));
    Odrv4 I__3141 (
            .O(N__17590),
            .I(\Lab_UT.dictrl.currState_ret_3and ));
    InMux I__3140 (
            .O(N__17587),
            .I(N__17584));
    LocalMux I__3139 (
            .O(N__17584),
            .I(N__17581));
    Span4Mux_h I__3138 (
            .O(N__17581),
            .I(N__17578));
    Span4Mux_h I__3137 (
            .O(N__17578),
            .I(N__17575));
    Odrv4 I__3136 (
            .O(N__17575),
            .I(\Lab_UT.dictrl.currState_0_ret_28_RNOZ0Z_2 ));
    InMux I__3135 (
            .O(N__17572),
            .I(N__17568));
    InMux I__3134 (
            .O(N__17571),
            .I(N__17562));
    LocalMux I__3133 (
            .O(N__17568),
            .I(N__17559));
    InMux I__3132 (
            .O(N__17567),
            .I(N__17554));
    InMux I__3131 (
            .O(N__17566),
            .I(N__17554));
    CascadeMux I__3130 (
            .O(N__17565),
            .I(N__17549));
    LocalMux I__3129 (
            .O(N__17562),
            .I(N__17543));
    Span4Mux_v I__3128 (
            .O(N__17559),
            .I(N__17538));
    LocalMux I__3127 (
            .O(N__17554),
            .I(N__17538));
    InMux I__3126 (
            .O(N__17553),
            .I(N__17533));
    InMux I__3125 (
            .O(N__17552),
            .I(N__17533));
    InMux I__3124 (
            .O(N__17549),
            .I(N__17527));
    InMux I__3123 (
            .O(N__17548),
            .I(N__17527));
    InMux I__3122 (
            .O(N__17547),
            .I(N__17521));
    InMux I__3121 (
            .O(N__17546),
            .I(N__17521));
    Span4Mux_h I__3120 (
            .O(N__17543),
            .I(N__17516));
    Span4Mux_h I__3119 (
            .O(N__17538),
            .I(N__17516));
    LocalMux I__3118 (
            .O(N__17533),
            .I(N__17513));
    InMux I__3117 (
            .O(N__17532),
            .I(N__17510));
    LocalMux I__3116 (
            .O(N__17527),
            .I(N__17507));
    InMux I__3115 (
            .O(N__17526),
            .I(N__17504));
    LocalMux I__3114 (
            .O(N__17521),
            .I(\Lab_UT.dictrl.N_8ctr ));
    Odrv4 I__3113 (
            .O(N__17516),
            .I(\Lab_UT.dictrl.N_8ctr ));
    Odrv4 I__3112 (
            .O(N__17513),
            .I(\Lab_UT.dictrl.N_8ctr ));
    LocalMux I__3111 (
            .O(N__17510),
            .I(\Lab_UT.dictrl.N_8ctr ));
    Odrv12 I__3110 (
            .O(N__17507),
            .I(\Lab_UT.dictrl.N_8ctr ));
    LocalMux I__3109 (
            .O(N__17504),
            .I(\Lab_UT.dictrl.N_8ctr ));
    CascadeMux I__3108 (
            .O(N__17491),
            .I(\Lab_UT.dictrl.currState_0_ret_28_RNOZ0Z_3_cascade_ ));
    InMux I__3107 (
            .O(N__17488),
            .I(N__17485));
    LocalMux I__3106 (
            .O(N__17485),
            .I(N__17482));
    Odrv4 I__3105 (
            .O(N__17482),
            .I(\Lab_UT.dictrl.N_8_0 ));
    InMux I__3104 (
            .O(N__17479),
            .I(N__17476));
    LocalMux I__3103 (
            .O(N__17476),
            .I(\Lab_UT.dictrl.r_dicLdMtens21_1_reti ));
    InMux I__3102 (
            .O(N__17473),
            .I(N__17469));
    InMux I__3101 (
            .O(N__17472),
            .I(N__17466));
    LocalMux I__3100 (
            .O(N__17469),
            .I(N__17461));
    LocalMux I__3099 (
            .O(N__17466),
            .I(N__17461));
    Odrv4 I__3098 (
            .O(N__17461),
            .I(\Lab_UT.dictrl.decoder.de_littleA_2Z0Z_0 ));
    CascadeMux I__3097 (
            .O(N__17458),
            .I(\Lab_UT.dictrl.de_littleA_1_cascade_ ));
    CascadeMux I__3096 (
            .O(N__17455),
            .I(\Lab_UT.dictrl.N_37_0_cascade_ ));
    InMux I__3095 (
            .O(N__17452),
            .I(N__17449));
    LocalMux I__3094 (
            .O(N__17449),
            .I(N__17446));
    Odrv4 I__3093 (
            .O(N__17446),
            .I(\Lab_UT.dictrl.g0_15_rn_1 ));
    InMux I__3092 (
            .O(N__17443),
            .I(N__17437));
    InMux I__3091 (
            .O(N__17442),
            .I(N__17437));
    LocalMux I__3090 (
            .O(N__17437),
            .I(N__17434));
    Span4Mux_h I__3089 (
            .O(N__17434),
            .I(N__17431));
    Odrv4 I__3088 (
            .O(N__17431),
            .I(\Lab_UT.dictrl.G_19_0_a7_0_1 ));
    InMux I__3087 (
            .O(N__17428),
            .I(N__17425));
    LocalMux I__3086 (
            .O(N__17425),
            .I(N__17422));
    Odrv12 I__3085 (
            .O(N__17422),
            .I(G_19_0_a7_4_7));
    InMux I__3084 (
            .O(N__17419),
            .I(N__17416));
    LocalMux I__3083 (
            .O(N__17416),
            .I(N__17412));
    InMux I__3082 (
            .O(N__17415),
            .I(N__17409));
    Odrv4 I__3081 (
            .O(N__17412),
            .I(\Lab_UT.dictrl.N_17_0 ));
    LocalMux I__3080 (
            .O(N__17409),
            .I(\Lab_UT.dictrl.N_17_0 ));
    CascadeMux I__3079 (
            .O(N__17404),
            .I(\Lab_UT.dictrl.N_13_cascade_ ));
    InMux I__3078 (
            .O(N__17401),
            .I(N__17398));
    LocalMux I__3077 (
            .O(N__17398),
            .I(N__17395));
    Span4Mux_v I__3076 (
            .O(N__17395),
            .I(N__17391));
    InMux I__3075 (
            .O(N__17394),
            .I(N__17388));
    Sp12to4 I__3074 (
            .O(N__17391),
            .I(N__17383));
    LocalMux I__3073 (
            .O(N__17388),
            .I(N__17383));
    Span12Mux_s10_h I__3072 (
            .O(N__17383),
            .I(N__17380));
    Odrv12 I__3071 (
            .O(N__17380),
            .I(\Lab_UT.dictrl.G_19_0_2 ));
    CascadeMux I__3070 (
            .O(N__17377),
            .I(\Lab_UT.dictrl.nextStateZ0Z_2_cascade_ ));
    InMux I__3069 (
            .O(N__17374),
            .I(N__17371));
    LocalMux I__3068 (
            .O(N__17371),
            .I(\Lab_UT.dictrl.dicLdASones_rst ));
    CascadeMux I__3067 (
            .O(N__17368),
            .I(\Lab_UT.dictrl.dicLdASones_rst_cascade_ ));
    InMux I__3066 (
            .O(N__17365),
            .I(N__17359));
    InMux I__3065 (
            .O(N__17364),
            .I(N__17359));
    LocalMux I__3064 (
            .O(N__17359),
            .I(\Lab_UT.dictrl.dicLdASonesZ0 ));
    CascadeMux I__3063 (
            .O(N__17356),
            .I(N__17352));
    InMux I__3062 (
            .O(N__17355),
            .I(N__17345));
    InMux I__3061 (
            .O(N__17352),
            .I(N__17345));
    InMux I__3060 (
            .O(N__17351),
            .I(N__17340));
    InMux I__3059 (
            .O(N__17350),
            .I(N__17340));
    LocalMux I__3058 (
            .O(N__17345),
            .I(\Lab_UT.dictrl.N_5ctr ));
    LocalMux I__3057 (
            .O(N__17340),
            .I(\Lab_UT.dictrl.N_5ctr ));
    CascadeMux I__3056 (
            .O(N__17335),
            .I(N__17332));
    InMux I__3055 (
            .O(N__17332),
            .I(N__17328));
    CascadeMux I__3054 (
            .O(N__17331),
            .I(N__17325));
    LocalMux I__3053 (
            .O(N__17328),
            .I(N__17322));
    InMux I__3052 (
            .O(N__17325),
            .I(N__17319));
    Span4Mux_v I__3051 (
            .O(N__17322),
            .I(N__17316));
    LocalMux I__3050 (
            .O(N__17319),
            .I(N__17313));
    Odrv4 I__3049 (
            .O(N__17316),
            .I(\Lab_UT.dictrl.N_7ctr ));
    Odrv4 I__3048 (
            .O(N__17313),
            .I(\Lab_UT.dictrl.N_7ctr ));
    InMux I__3047 (
            .O(N__17308),
            .I(N__17293));
    InMux I__3046 (
            .O(N__17307),
            .I(N__17293));
    InMux I__3045 (
            .O(N__17306),
            .I(N__17293));
    InMux I__3044 (
            .O(N__17305),
            .I(N__17293));
    InMux I__3043 (
            .O(N__17304),
            .I(N__17290));
    InMux I__3042 (
            .O(N__17303),
            .I(N__17285));
    InMux I__3041 (
            .O(N__17302),
            .I(N__17285));
    LocalMux I__3040 (
            .O(N__17293),
            .I(N__17282));
    LocalMux I__3039 (
            .O(N__17290),
            .I(N__17277));
    LocalMux I__3038 (
            .O(N__17285),
            .I(N__17277));
    Span4Mux_v I__3037 (
            .O(N__17282),
            .I(N__17274));
    Span4Mux_h I__3036 (
            .O(N__17277),
            .I(N__17271));
    Odrv4 I__3035 (
            .O(N__17274),
            .I(\Lab_UT.dictrl.nextState_RNIGHD18Z0Z_1 ));
    Odrv4 I__3034 (
            .O(N__17271),
            .I(\Lab_UT.dictrl.nextState_RNIGHD18Z0Z_1 ));
    InMux I__3033 (
            .O(N__17266),
            .I(N__17254));
    InMux I__3032 (
            .O(N__17265),
            .I(N__17247));
    InMux I__3031 (
            .O(N__17264),
            .I(N__17247));
    InMux I__3030 (
            .O(N__17263),
            .I(N__17247));
    InMux I__3029 (
            .O(N__17262),
            .I(N__17244));
    InMux I__3028 (
            .O(N__17261),
            .I(N__17241));
    InMux I__3027 (
            .O(N__17260),
            .I(N__17232));
    InMux I__3026 (
            .O(N__17259),
            .I(N__17232));
    InMux I__3025 (
            .O(N__17258),
            .I(N__17232));
    InMux I__3024 (
            .O(N__17257),
            .I(N__17232));
    LocalMux I__3023 (
            .O(N__17254),
            .I(N__17225));
    LocalMux I__3022 (
            .O(N__17247),
            .I(N__17225));
    LocalMux I__3021 (
            .O(N__17244),
            .I(N__17222));
    LocalMux I__3020 (
            .O(N__17241),
            .I(N__17216));
    LocalMux I__3019 (
            .O(N__17232),
            .I(N__17216));
    InMux I__3018 (
            .O(N__17231),
            .I(N__17213));
    InMux I__3017 (
            .O(N__17230),
            .I(N__17210));
    Span4Mux_h I__3016 (
            .O(N__17225),
            .I(N__17205));
    Span4Mux_s3_h I__3015 (
            .O(N__17222),
            .I(N__17205));
    InMux I__3014 (
            .O(N__17221),
            .I(N__17202));
    Span4Mux_s3_h I__3013 (
            .O(N__17216),
            .I(N__17199));
    LocalMux I__3012 (
            .O(N__17213),
            .I(N__17194));
    LocalMux I__3011 (
            .O(N__17210),
            .I(N__17194));
    Odrv4 I__3010 (
            .O(N__17205),
            .I(\Lab_UT.dictrl.i8_mux ));
    LocalMux I__3009 (
            .O(N__17202),
            .I(\Lab_UT.dictrl.i8_mux ));
    Odrv4 I__3008 (
            .O(N__17199),
            .I(\Lab_UT.dictrl.i8_mux ));
    Odrv12 I__3007 (
            .O(N__17194),
            .I(\Lab_UT.dictrl.i8_mux ));
    CascadeMux I__3006 (
            .O(N__17185),
            .I(N__17178));
    CascadeMux I__3005 (
            .O(N__17184),
            .I(N__17175));
    CascadeMux I__3004 (
            .O(N__17183),
            .I(N__17172));
    CascadeMux I__3003 (
            .O(N__17182),
            .I(N__17169));
    CascadeMux I__3002 (
            .O(N__17181),
            .I(N__17166));
    InMux I__3001 (
            .O(N__17178),
            .I(N__17161));
    InMux I__3000 (
            .O(N__17175),
            .I(N__17161));
    InMux I__2999 (
            .O(N__17172),
            .I(N__17156));
    InMux I__2998 (
            .O(N__17169),
            .I(N__17156));
    InMux I__2997 (
            .O(N__17166),
            .I(N__17153));
    LocalMux I__2996 (
            .O(N__17161),
            .I(N__17148));
    LocalMux I__2995 (
            .O(N__17156),
            .I(N__17148));
    LocalMux I__2994 (
            .O(N__17153),
            .I(N__17145));
    Span4Mux_h I__2993 (
            .O(N__17148),
            .I(N__17142));
    Odrv12 I__2992 (
            .O(N__17145),
            .I(\Lab_UT.dictrl.currState_2_RNI1O2A_0Z0Z_1 ));
    Odrv4 I__2991 (
            .O(N__17142),
            .I(\Lab_UT.dictrl.currState_2_RNI1O2A_0Z0Z_1 ));
    InMux I__2990 (
            .O(N__17137),
            .I(N__17134));
    LocalMux I__2989 (
            .O(N__17134),
            .I(N__17131));
    Odrv12 I__2988 (
            .O(N__17131),
            .I(\Lab_UT.dictrl.g0_13_1 ));
    InMux I__2987 (
            .O(N__17128),
            .I(N__17125));
    LocalMux I__2986 (
            .O(N__17125),
            .I(\Lab_UT.dictrl.g0_1 ));
    InMux I__2985 (
            .O(N__17122),
            .I(N__17119));
    LocalMux I__2984 (
            .O(N__17119),
            .I(\Lab_UT.dictrl.g0_i_o4_0_0 ));
    CascadeMux I__2983 (
            .O(N__17116),
            .I(\Lab_UT.dictrl.currState_0_ret_20and_1_0_cascade_ ));
    InMux I__2982 (
            .O(N__17113),
            .I(N__17109));
    InMux I__2981 (
            .O(N__17112),
            .I(N__17106));
    LocalMux I__2980 (
            .O(N__17109),
            .I(N__17103));
    LocalMux I__2979 (
            .O(N__17106),
            .I(N__17100));
    Span4Mux_v I__2978 (
            .O(N__17103),
            .I(N__17094));
    Span4Mux_s2_h I__2977 (
            .O(N__17100),
            .I(N__17094));
    InMux I__2976 (
            .O(N__17099),
            .I(N__17091));
    Span4Mux_h I__2975 (
            .O(N__17094),
            .I(N__17088));
    LocalMux I__2974 (
            .O(N__17091),
            .I(\Lab_UT.dictrl.de_cr ));
    Odrv4 I__2973 (
            .O(N__17088),
            .I(\Lab_UT.dictrl.de_cr ));
    CascadeMux I__2972 (
            .O(N__17083),
            .I(N__17080));
    InMux I__2971 (
            .O(N__17080),
            .I(N__17077));
    LocalMux I__2970 (
            .O(N__17077),
            .I(N__17074));
    Odrv4 I__2969 (
            .O(N__17074),
            .I(\Lab_UT.dictrl.N_13 ));
    CascadeMux I__2968 (
            .O(N__17071),
            .I(N__17068));
    InMux I__2967 (
            .O(N__17068),
            .I(N__17065));
    LocalMux I__2966 (
            .O(N__17065),
            .I(N__17062));
    Span4Mux_h I__2965 (
            .O(N__17062),
            .I(N__17059));
    Odrv4 I__2964 (
            .O(N__17059),
            .I(\Lab_UT.N_91 ));
    InMux I__2963 (
            .O(N__17056),
            .I(N__17053));
    LocalMux I__2962 (
            .O(N__17053),
            .I(N__17050));
    Span4Mux_h I__2961 (
            .O(N__17050),
            .I(N__17047));
    Odrv4 I__2960 (
            .O(N__17047),
            .I(\Lab_UT.N_83 ));
    CascadeMux I__2959 (
            .O(N__17044),
            .I(N__17034));
    InMux I__2958 (
            .O(N__17043),
            .I(N__17023));
    InMux I__2957 (
            .O(N__17042),
            .I(N__17023));
    InMux I__2956 (
            .O(N__17041),
            .I(N__17023));
    InMux I__2955 (
            .O(N__17040),
            .I(N__17023));
    InMux I__2954 (
            .O(N__17039),
            .I(N__17012));
    InMux I__2953 (
            .O(N__17038),
            .I(N__17012));
    InMux I__2952 (
            .O(N__17037),
            .I(N__17012));
    InMux I__2951 (
            .O(N__17034),
            .I(N__17012));
    InMux I__2950 (
            .O(N__17033),
            .I(N__17012));
    InMux I__2949 (
            .O(N__17032),
            .I(N__17009));
    LocalMux I__2948 (
            .O(N__17023),
            .I(\Lab_UT.Mten_at_0 ));
    LocalMux I__2947 (
            .O(N__17012),
            .I(\Lab_UT.Mten_at_0 ));
    LocalMux I__2946 (
            .O(N__17009),
            .I(\Lab_UT.Mten_at_0 ));
    CascadeMux I__2945 (
            .O(N__17002),
            .I(N__16995));
    CascadeMux I__2944 (
            .O(N__17001),
            .I(N__16991));
    CascadeMux I__2943 (
            .O(N__17000),
            .I(N__16988));
    CascadeMux I__2942 (
            .O(N__16999),
            .I(N__16984));
    CascadeMux I__2941 (
            .O(N__16998),
            .I(N__16980));
    InMux I__2940 (
            .O(N__16995),
            .I(N__16970));
    InMux I__2939 (
            .O(N__16994),
            .I(N__16970));
    InMux I__2938 (
            .O(N__16991),
            .I(N__16970));
    InMux I__2937 (
            .O(N__16988),
            .I(N__16970));
    InMux I__2936 (
            .O(N__16987),
            .I(N__16967));
    InMux I__2935 (
            .O(N__16984),
            .I(N__16958));
    InMux I__2934 (
            .O(N__16983),
            .I(N__16958));
    InMux I__2933 (
            .O(N__16980),
            .I(N__16958));
    InMux I__2932 (
            .O(N__16979),
            .I(N__16958));
    LocalMux I__2931 (
            .O(N__16970),
            .I(\Lab_UT.Mten_at_3 ));
    LocalMux I__2930 (
            .O(N__16967),
            .I(\Lab_UT.Mten_at_3 ));
    LocalMux I__2929 (
            .O(N__16958),
            .I(\Lab_UT.Mten_at_3 ));
    CascadeMux I__2928 (
            .O(N__16951),
            .I(\Lab_UT.Mten_at_0_cascade_ ));
    InMux I__2927 (
            .O(N__16948),
            .I(N__16945));
    LocalMux I__2926 (
            .O(N__16945),
            .I(\Lab_UT.N_77 ));
    InMux I__2925 (
            .O(N__16942),
            .I(N__16925));
    InMux I__2924 (
            .O(N__16941),
            .I(N__16925));
    InMux I__2923 (
            .O(N__16940),
            .I(N__16925));
    InMux I__2922 (
            .O(N__16939),
            .I(N__16925));
    InMux I__2921 (
            .O(N__16938),
            .I(N__16922));
    InMux I__2920 (
            .O(N__16937),
            .I(N__16913));
    InMux I__2919 (
            .O(N__16936),
            .I(N__16913));
    InMux I__2918 (
            .O(N__16935),
            .I(N__16913));
    InMux I__2917 (
            .O(N__16934),
            .I(N__16913));
    LocalMux I__2916 (
            .O(N__16925),
            .I(\Lab_UT.Mten_at_1 ));
    LocalMux I__2915 (
            .O(N__16922),
            .I(\Lab_UT.Mten_at_1 ));
    LocalMux I__2914 (
            .O(N__16913),
            .I(\Lab_UT.Mten_at_1 ));
    InMux I__2913 (
            .O(N__16906),
            .I(N__16903));
    LocalMux I__2912 (
            .O(N__16903),
            .I(\Lab_UT.N_77_1 ));
    InMux I__2911 (
            .O(N__16900),
            .I(N__16897));
    LocalMux I__2910 (
            .O(N__16897),
            .I(\uu2.bitmapZ0Z_84 ));
    InMux I__2909 (
            .O(N__16894),
            .I(N__16891));
    LocalMux I__2908 (
            .O(N__16891),
            .I(N__16888));
    Span4Mux_h I__2907 (
            .O(N__16888),
            .I(N__16885));
    Odrv4 I__2906 (
            .O(N__16885),
            .I(\Lab_UT.L3_segment4_0_i_1_5 ));
    InMux I__2905 (
            .O(N__16882),
            .I(N__16879));
    LocalMux I__2904 (
            .O(N__16879),
            .I(N__16876));
    Odrv4 I__2903 (
            .O(N__16876),
            .I(\Lab_UT.N_65 ));
    CascadeMux I__2902 (
            .O(N__16873),
            .I(\Lab_UT.Mten_at_3_cascade_ ));
    InMux I__2901 (
            .O(N__16870),
            .I(N__16867));
    LocalMux I__2900 (
            .O(N__16867),
            .I(N__16864));
    Span4Mux_h I__2899 (
            .O(N__16864),
            .I(N__16861));
    Odrv4 I__2898 (
            .O(N__16861),
            .I(\Lab_UT.segment_1_3 ));
    InMux I__2897 (
            .O(N__16858),
            .I(N__16852));
    InMux I__2896 (
            .O(N__16857),
            .I(N__16852));
    LocalMux I__2895 (
            .O(N__16852),
            .I(\Lab_UT.N_69_0 ));
    CascadeMux I__2894 (
            .O(N__16849),
            .I(\Lab_UT.N_69_0_cascade_ ));
    InMux I__2893 (
            .O(N__16846),
            .I(N__16843));
    LocalMux I__2892 (
            .O(N__16843),
            .I(N__16840));
    Span4Mux_h I__2891 (
            .O(N__16840),
            .I(N__16837));
    Odrv4 I__2890 (
            .O(N__16837),
            .I(\Lab_UT.N_92 ));
    InMux I__2889 (
            .O(N__16834),
            .I(N__16828));
    InMux I__2888 (
            .O(N__16833),
            .I(N__16828));
    LocalMux I__2887 (
            .O(N__16828),
            .I(\Lab_UT.N_67_0 ));
    CascadeMux I__2886 (
            .O(N__16825),
            .I(\Lab_UT.N_65_2_cascade_ ));
    InMux I__2885 (
            .O(N__16822),
            .I(N__16819));
    LocalMux I__2884 (
            .O(N__16819),
            .I(\Lab_UT.segment_1_2_6 ));
    InMux I__2883 (
            .O(N__16816),
            .I(N__16813));
    LocalMux I__2882 (
            .O(N__16813),
            .I(N__16810));
    Odrv4 I__2881 (
            .O(N__16810),
            .I(\uu2.bitmapZ0Z_186 ));
    CascadeMux I__2880 (
            .O(N__16807),
            .I(\Lab_UT.N_76_2_cascade_ ));
    InMux I__2879 (
            .O(N__16804),
            .I(N__16801));
    LocalMux I__2878 (
            .O(N__16801),
            .I(\uu2.bitmapZ0Z_90 ));
    CascadeMux I__2877 (
            .O(N__16798),
            .I(N__16795));
    InMux I__2876 (
            .O(N__16795),
            .I(N__16792));
    LocalMux I__2875 (
            .O(N__16792),
            .I(\uu2.bitmapZ0Z_218 ));
    InMux I__2874 (
            .O(N__16789),
            .I(N__16781));
    InMux I__2873 (
            .O(N__16788),
            .I(N__16781));
    InMux I__2872 (
            .O(N__16787),
            .I(N__16772));
    InMux I__2871 (
            .O(N__16786),
            .I(N__16772));
    LocalMux I__2870 (
            .O(N__16781),
            .I(N__16764));
    InMux I__2869 (
            .O(N__16780),
            .I(N__16761));
    CascadeMux I__2868 (
            .O(N__16779),
            .I(N__16758));
    InMux I__2867 (
            .O(N__16778),
            .I(N__16751));
    InMux I__2866 (
            .O(N__16777),
            .I(N__16751));
    LocalMux I__2865 (
            .O(N__16772),
            .I(N__16748));
    InMux I__2864 (
            .O(N__16771),
            .I(N__16745));
    InMux I__2863 (
            .O(N__16770),
            .I(N__16740));
    InMux I__2862 (
            .O(N__16769),
            .I(N__16740));
    InMux I__2861 (
            .O(N__16768),
            .I(N__16737));
    InMux I__2860 (
            .O(N__16767),
            .I(N__16734));
    Span4Mux_h I__2859 (
            .O(N__16764),
            .I(N__16731));
    LocalMux I__2858 (
            .O(N__16761),
            .I(N__16728));
    InMux I__2857 (
            .O(N__16758),
            .I(N__16721));
    InMux I__2856 (
            .O(N__16757),
            .I(N__16721));
    InMux I__2855 (
            .O(N__16756),
            .I(N__16721));
    LocalMux I__2854 (
            .O(N__16751),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    Odrv4 I__2853 (
            .O(N__16748),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    LocalMux I__2852 (
            .O(N__16745),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    LocalMux I__2851 (
            .O(N__16740),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    LocalMux I__2850 (
            .O(N__16737),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    LocalMux I__2849 (
            .O(N__16734),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    Odrv4 I__2848 (
            .O(N__16731),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    Odrv4 I__2847 (
            .O(N__16728),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    LocalMux I__2846 (
            .O(N__16721),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    CascadeMux I__2845 (
            .O(N__16702),
            .I(\Lab_UT.N_76_1_cascade_ ));
    InMux I__2844 (
            .O(N__16699),
            .I(N__16696));
    LocalMux I__2843 (
            .O(N__16696),
            .I(N__16693));
    Span4Mux_h I__2842 (
            .O(N__16693),
            .I(N__16690));
    Odrv4 I__2841 (
            .O(N__16690),
            .I(\uu2.bitmapZ0Z_212 ));
    CascadeMux I__2840 (
            .O(N__16687),
            .I(\Lab_UT.N_65_1_cascade_ ));
    InMux I__2839 (
            .O(N__16684),
            .I(N__16681));
    LocalMux I__2838 (
            .O(N__16681),
            .I(\Lab_UT.segment_1_1_6 ));
    InMux I__2837 (
            .O(N__16678),
            .I(N__16675));
    LocalMux I__2836 (
            .O(N__16675),
            .I(\uu2.bitmapZ0Z_180 ));
    CascadeMux I__2835 (
            .O(N__16672),
            .I(\Lab_UT.L3_segment2_1_2_cascade_ ));
    CascadeMux I__2834 (
            .O(N__16669),
            .I(N__16666));
    InMux I__2833 (
            .O(N__16666),
            .I(N__16663));
    LocalMux I__2832 (
            .O(N__16663),
            .I(N__16660));
    Span4Mux_v I__2831 (
            .O(N__16660),
            .I(N__16657));
    Odrv4 I__2830 (
            .O(N__16657),
            .I(\uu2.bitmapZ0Z_215 ));
    CascadeMux I__2829 (
            .O(N__16654),
            .I(\Lab_UT.L3_segment2_0_i_1_0_cascade_ ));
    InMux I__2828 (
            .O(N__16651),
            .I(N__16648));
    LocalMux I__2827 (
            .O(N__16648),
            .I(\uu2.bitmapZ0Z_52 ));
    InMux I__2826 (
            .O(N__16645),
            .I(N__16636));
    InMux I__2825 (
            .O(N__16644),
            .I(N__16633));
    InMux I__2824 (
            .O(N__16643),
            .I(N__16628));
    InMux I__2823 (
            .O(N__16642),
            .I(N__16628));
    InMux I__2822 (
            .O(N__16641),
            .I(N__16622));
    InMux I__2821 (
            .O(N__16640),
            .I(N__16622));
    CascadeMux I__2820 (
            .O(N__16639),
            .I(N__16619));
    LocalMux I__2819 (
            .O(N__16636),
            .I(N__16613));
    LocalMux I__2818 (
            .O(N__16633),
            .I(N__16608));
    LocalMux I__2817 (
            .O(N__16628),
            .I(N__16608));
    InMux I__2816 (
            .O(N__16627),
            .I(N__16605));
    LocalMux I__2815 (
            .O(N__16622),
            .I(N__16601));
    InMux I__2814 (
            .O(N__16619),
            .I(N__16598));
    InMux I__2813 (
            .O(N__16618),
            .I(N__16595));
    InMux I__2812 (
            .O(N__16617),
            .I(N__16590));
    InMux I__2811 (
            .O(N__16616),
            .I(N__16590));
    Span4Mux_s3_v I__2810 (
            .O(N__16613),
            .I(N__16583));
    Span4Mux_v I__2809 (
            .O(N__16608),
            .I(N__16583));
    LocalMux I__2808 (
            .O(N__16605),
            .I(N__16583));
    InMux I__2807 (
            .O(N__16604),
            .I(N__16580));
    Span4Mux_h I__2806 (
            .O(N__16601),
            .I(N__16577));
    LocalMux I__2805 (
            .O(N__16598),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    LocalMux I__2804 (
            .O(N__16595),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    LocalMux I__2803 (
            .O(N__16590),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    Odrv4 I__2802 (
            .O(N__16583),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    LocalMux I__2801 (
            .O(N__16580),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    Odrv4 I__2800 (
            .O(N__16577),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    InMux I__2799 (
            .O(N__16564),
            .I(N__16561));
    LocalMux I__2798 (
            .O(N__16561),
            .I(\uu2.bitmapZ0Z_308 ));
    InMux I__2797 (
            .O(N__16558),
            .I(N__16555));
    LocalMux I__2796 (
            .O(N__16555),
            .I(\uu2.N_158 ));
    CascadeMux I__2795 (
            .O(N__16552),
            .I(\Lab_UT.segmentUQ_0_0_1_cascade_ ));
    InMux I__2794 (
            .O(N__16549),
            .I(N__16546));
    LocalMux I__2793 (
            .O(N__16546),
            .I(N__16540));
    InMux I__2792 (
            .O(N__16545),
            .I(N__16537));
    CascadeMux I__2791 (
            .O(N__16544),
            .I(N__16534));
    InMux I__2790 (
            .O(N__16543),
            .I(N__16530));
    Span4Mux_v I__2789 (
            .O(N__16540),
            .I(N__16525));
    LocalMux I__2788 (
            .O(N__16537),
            .I(N__16525));
    InMux I__2787 (
            .O(N__16534),
            .I(N__16520));
    InMux I__2786 (
            .O(N__16533),
            .I(N__16520));
    LocalMux I__2785 (
            .O(N__16530),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    Odrv4 I__2784 (
            .O(N__16525),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    LocalMux I__2783 (
            .O(N__16520),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    InMux I__2782 (
            .O(N__16513),
            .I(N__16507));
    InMux I__2781 (
            .O(N__16512),
            .I(N__16507));
    LocalMux I__2780 (
            .O(N__16507),
            .I(N__16501));
    InMux I__2779 (
            .O(N__16506),
            .I(N__16495));
    InMux I__2778 (
            .O(N__16505),
            .I(N__16492));
    InMux I__2777 (
            .O(N__16504),
            .I(N__16489));
    Span4Mux_h I__2776 (
            .O(N__16501),
            .I(N__16486));
    InMux I__2775 (
            .O(N__16500),
            .I(N__16481));
    InMux I__2774 (
            .O(N__16499),
            .I(N__16481));
    InMux I__2773 (
            .O(N__16498),
            .I(N__16478));
    LocalMux I__2772 (
            .O(N__16495),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    LocalMux I__2771 (
            .O(N__16492),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    LocalMux I__2770 (
            .O(N__16489),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    Odrv4 I__2769 (
            .O(N__16486),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    LocalMux I__2768 (
            .O(N__16481),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    LocalMux I__2767 (
            .O(N__16478),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    InMux I__2766 (
            .O(N__16465),
            .I(N__16462));
    LocalMux I__2765 (
            .O(N__16462),
            .I(N__16458));
    InMux I__2764 (
            .O(N__16461),
            .I(N__16455));
    Span4Mux_v I__2763 (
            .O(N__16458),
            .I(N__16452));
    LocalMux I__2762 (
            .O(N__16455),
            .I(\uu2.N_41 ));
    Odrv4 I__2761 (
            .O(N__16452),
            .I(\uu2.N_41 ));
    CascadeMux I__2760 (
            .O(N__16447),
            .I(N__16443));
    InMux I__2759 (
            .O(N__16446),
            .I(N__16437));
    InMux I__2758 (
            .O(N__16443),
            .I(N__16434));
    CascadeMux I__2757 (
            .O(N__16442),
            .I(N__16430));
    InMux I__2756 (
            .O(N__16441),
            .I(N__16425));
    InMux I__2755 (
            .O(N__16440),
            .I(N__16425));
    LocalMux I__2754 (
            .O(N__16437),
            .I(N__16422));
    LocalMux I__2753 (
            .O(N__16434),
            .I(N__16419));
    InMux I__2752 (
            .O(N__16433),
            .I(N__16416));
    InMux I__2751 (
            .O(N__16430),
            .I(N__16413));
    LocalMux I__2750 (
            .O(N__16425),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    Odrv4 I__2749 (
            .O(N__16422),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    Odrv4 I__2748 (
            .O(N__16419),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    LocalMux I__2747 (
            .O(N__16416),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    LocalMux I__2746 (
            .O(N__16413),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    CascadeMux I__2745 (
            .O(N__16402),
            .I(\uu2.N_41_cascade_ ));
    InMux I__2744 (
            .O(N__16399),
            .I(N__16392));
    InMux I__2743 (
            .O(N__16398),
            .I(N__16392));
    CascadeMux I__2742 (
            .O(N__16397),
            .I(N__16389));
    LocalMux I__2741 (
            .O(N__16392),
            .I(N__16385));
    InMux I__2740 (
            .O(N__16389),
            .I(N__16380));
    InMux I__2739 (
            .O(N__16388),
            .I(N__16380));
    Odrv4 I__2738 (
            .O(N__16385),
            .I(\uu2.N_43 ));
    LocalMux I__2737 (
            .O(N__16380),
            .I(\uu2.N_43 ));
    InMux I__2736 (
            .O(N__16375),
            .I(N__16371));
    CascadeMux I__2735 (
            .O(N__16374),
            .I(N__16368));
    LocalMux I__2734 (
            .O(N__16371),
            .I(N__16365));
    InMux I__2733 (
            .O(N__16368),
            .I(N__16358));
    Span4Mux_v I__2732 (
            .O(N__16365),
            .I(N__16355));
    InMux I__2731 (
            .O(N__16364),
            .I(N__16346));
    InMux I__2730 (
            .O(N__16363),
            .I(N__16346));
    InMux I__2729 (
            .O(N__16362),
            .I(N__16346));
    InMux I__2728 (
            .O(N__16361),
            .I(N__16346));
    LocalMux I__2727 (
            .O(N__16358),
            .I(\uu2.N_40 ));
    Odrv4 I__2726 (
            .O(N__16355),
            .I(\uu2.N_40 ));
    LocalMux I__2725 (
            .O(N__16346),
            .I(\uu2.N_40 ));
    CascadeMux I__2724 (
            .O(N__16339),
            .I(\uu2.N_43_cascade_ ));
    CascadeMux I__2723 (
            .O(N__16336),
            .I(N__16333));
    InMux I__2722 (
            .O(N__16333),
            .I(N__16326));
    InMux I__2721 (
            .O(N__16332),
            .I(N__16323));
    InMux I__2720 (
            .O(N__16331),
            .I(N__16316));
    InMux I__2719 (
            .O(N__16330),
            .I(N__16316));
    InMux I__2718 (
            .O(N__16329),
            .I(N__16316));
    LocalMux I__2717 (
            .O(N__16326),
            .I(N__16311));
    LocalMux I__2716 (
            .O(N__16323),
            .I(N__16311));
    LocalMux I__2715 (
            .O(N__16316),
            .I(\uu2.w_addr_displaying_RNIFCPV4Z0Z_8 ));
    Odrv4 I__2714 (
            .O(N__16311),
            .I(\uu2.w_addr_displaying_RNIFCPV4Z0Z_8 ));
    CascadeMux I__2713 (
            .O(N__16306),
            .I(\uu2.w_addr_displaying_RNIFCPV4Z0Z_8_cascade_ ));
    CEMux I__2712 (
            .O(N__16303),
            .I(N__16300));
    LocalMux I__2711 (
            .O(N__16300),
            .I(N__16297));
    Odrv4 I__2710 (
            .O(N__16297),
            .I(\uu2.N_36_0 ));
    InMux I__2709 (
            .O(N__16294),
            .I(N__16291));
    LocalMux I__2708 (
            .O(N__16291),
            .I(\Lab_UT.L3_segment2_1_1 ));
    CascadeMux I__2707 (
            .O(N__16288),
            .I(\Lab_UT.L3_segment2_0_i_1_3_cascade_ ));
    CascadeMux I__2706 (
            .O(N__16285),
            .I(\uu2.un3_w_addr_user_4_cascade_ ));
    InMux I__2705 (
            .O(N__16282),
            .I(N__16279));
    LocalMux I__2704 (
            .O(N__16279),
            .I(\uu2.un3_w_addr_user_5 ));
    InMux I__2703 (
            .O(N__16276),
            .I(N__16268));
    InMux I__2702 (
            .O(N__16275),
            .I(N__16260));
    InMux I__2701 (
            .O(N__16274),
            .I(N__16260));
    InMux I__2700 (
            .O(N__16273),
            .I(N__16260));
    CascadeMux I__2699 (
            .O(N__16272),
            .I(N__16247));
    InMux I__2698 (
            .O(N__16271),
            .I(N__16244));
    LocalMux I__2697 (
            .O(N__16268),
            .I(N__16241));
    InMux I__2696 (
            .O(N__16267),
            .I(N__16238));
    LocalMux I__2695 (
            .O(N__16260),
            .I(N__16235));
    InMux I__2694 (
            .O(N__16259),
            .I(N__16232));
    InMux I__2693 (
            .O(N__16258),
            .I(N__16227));
    InMux I__2692 (
            .O(N__16257),
            .I(N__16227));
    InMux I__2691 (
            .O(N__16256),
            .I(N__16218));
    InMux I__2690 (
            .O(N__16255),
            .I(N__16218));
    InMux I__2689 (
            .O(N__16254),
            .I(N__16218));
    InMux I__2688 (
            .O(N__16253),
            .I(N__16218));
    InMux I__2687 (
            .O(N__16252),
            .I(N__16209));
    InMux I__2686 (
            .O(N__16251),
            .I(N__16209));
    InMux I__2685 (
            .O(N__16250),
            .I(N__16209));
    InMux I__2684 (
            .O(N__16247),
            .I(N__16209));
    LocalMux I__2683 (
            .O(N__16244),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    Odrv4 I__2682 (
            .O(N__16241),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    LocalMux I__2681 (
            .O(N__16238),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    Odrv4 I__2680 (
            .O(N__16235),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    LocalMux I__2679 (
            .O(N__16232),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    LocalMux I__2678 (
            .O(N__16227),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    LocalMux I__2677 (
            .O(N__16218),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    LocalMux I__2676 (
            .O(N__16209),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    CascadeMux I__2675 (
            .O(N__16192),
            .I(N__16189));
    InMux I__2674 (
            .O(N__16189),
            .I(N__16186));
    LocalMux I__2673 (
            .O(N__16186),
            .I(N__16183));
    Odrv12 I__2672 (
            .O(N__16183),
            .I(\uu2.mem0.w_addr_3 ));
    CascadeMux I__2671 (
            .O(N__16180),
            .I(\uu2.vbuf_w_addr_user.un448_ci_0_cascade_ ));
    InMux I__2670 (
            .O(N__16177),
            .I(N__16174));
    LocalMux I__2669 (
            .O(N__16174),
            .I(N__16169));
    InMux I__2668 (
            .O(N__16173),
            .I(N__16164));
    InMux I__2667 (
            .O(N__16172),
            .I(N__16164));
    Odrv4 I__2666 (
            .O(N__16169),
            .I(\uu2.w_addr_userZ0Z_8 ));
    LocalMux I__2665 (
            .O(N__16164),
            .I(\uu2.w_addr_userZ0Z_8 ));
    InMux I__2664 (
            .O(N__16159),
            .I(N__16156));
    LocalMux I__2663 (
            .O(N__16156),
            .I(N__16152));
    CascadeMux I__2662 (
            .O(N__16155),
            .I(N__16147));
    Span4Mux_h I__2661 (
            .O(N__16152),
            .I(N__16144));
    InMux I__2660 (
            .O(N__16151),
            .I(N__16137));
    InMux I__2659 (
            .O(N__16150),
            .I(N__16137));
    InMux I__2658 (
            .O(N__16147),
            .I(N__16137));
    Odrv4 I__2657 (
            .O(N__16144),
            .I(\uu2.w_addr_userZ0Z_7 ));
    LocalMux I__2656 (
            .O(N__16137),
            .I(\uu2.w_addr_userZ0Z_7 ));
    InMux I__2655 (
            .O(N__16132),
            .I(N__16122));
    InMux I__2654 (
            .O(N__16131),
            .I(N__16122));
    InMux I__2653 (
            .O(N__16130),
            .I(N__16122));
    InMux I__2652 (
            .O(N__16129),
            .I(N__16115));
    LocalMux I__2651 (
            .O(N__16122),
            .I(N__16112));
    CascadeMux I__2650 (
            .O(N__16121),
            .I(N__16105));
    InMux I__2649 (
            .O(N__16120),
            .I(N__16098));
    InMux I__2648 (
            .O(N__16119),
            .I(N__16098));
    InMux I__2647 (
            .O(N__16118),
            .I(N__16095));
    LocalMux I__2646 (
            .O(N__16115),
            .I(N__16092));
    Span4Mux_h I__2645 (
            .O(N__16112),
            .I(N__16089));
    InMux I__2644 (
            .O(N__16111),
            .I(N__16084));
    InMux I__2643 (
            .O(N__16110),
            .I(N__16084));
    InMux I__2642 (
            .O(N__16109),
            .I(N__16081));
    InMux I__2641 (
            .O(N__16108),
            .I(N__16072));
    InMux I__2640 (
            .O(N__16105),
            .I(N__16072));
    InMux I__2639 (
            .O(N__16104),
            .I(N__16072));
    InMux I__2638 (
            .O(N__16103),
            .I(N__16072));
    LocalMux I__2637 (
            .O(N__16098),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    LocalMux I__2636 (
            .O(N__16095),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    Odrv4 I__2635 (
            .O(N__16092),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    Odrv4 I__2634 (
            .O(N__16089),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    LocalMux I__2633 (
            .O(N__16084),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    LocalMux I__2632 (
            .O(N__16081),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    LocalMux I__2631 (
            .O(N__16072),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    CascadeMux I__2630 (
            .O(N__16057),
            .I(N__16054));
    InMux I__2629 (
            .O(N__16054),
            .I(N__16047));
    InMux I__2628 (
            .O(N__16053),
            .I(N__16047));
    CascadeMux I__2627 (
            .O(N__16052),
            .I(N__16044));
    LocalMux I__2626 (
            .O(N__16047),
            .I(N__16041));
    InMux I__2625 (
            .O(N__16044),
            .I(N__16038));
    Odrv4 I__2624 (
            .O(N__16041),
            .I(\uu2.N_39 ));
    LocalMux I__2623 (
            .O(N__16038),
            .I(\uu2.N_39 ));
    InMux I__2622 (
            .O(N__16033),
            .I(N__16030));
    LocalMux I__2621 (
            .O(N__16030),
            .I(N__16026));
    InMux I__2620 (
            .O(N__16029),
            .I(N__16023));
    Span4Mux_h I__2619 (
            .O(N__16026),
            .I(N__16020));
    LocalMux I__2618 (
            .O(N__16023),
            .I(\Lab_UT.uu0.l_countZ0Z_13 ));
    Odrv4 I__2617 (
            .O(N__16020),
            .I(\Lab_UT.uu0.l_countZ0Z_13 ));
    CascadeMux I__2616 (
            .O(N__16015),
            .I(\Lab_UT.uu0.un143_ci_0_cascade_ ));
    CascadeMux I__2615 (
            .O(N__16012),
            .I(\Lab_UT.uu0.un154_ci_9_cascade_ ));
    InMux I__2614 (
            .O(N__16009),
            .I(N__16006));
    LocalMux I__2613 (
            .O(N__16006),
            .I(N__16001));
    InMux I__2612 (
            .O(N__16005),
            .I(N__15996));
    InMux I__2611 (
            .O(N__16004),
            .I(N__15996));
    Span4Mux_h I__2610 (
            .O(N__16001),
            .I(N__15993));
    LocalMux I__2609 (
            .O(N__15996),
            .I(\Lab_UT.uu0.l_countZ0Z_12 ));
    Odrv4 I__2608 (
            .O(N__15993),
            .I(\Lab_UT.uu0.l_countZ0Z_12 ));
    CascadeMux I__2607 (
            .O(N__15988),
            .I(N__15985));
    InMux I__2606 (
            .O(N__15985),
            .I(N__15982));
    LocalMux I__2605 (
            .O(N__15982),
            .I(\Lab_UT.uu0.un165_ci_0 ));
    InMux I__2604 (
            .O(N__15979),
            .I(N__15955));
    InMux I__2603 (
            .O(N__15978),
            .I(N__15955));
    InMux I__2602 (
            .O(N__15977),
            .I(N__15955));
    InMux I__2601 (
            .O(N__15976),
            .I(N__15955));
    InMux I__2600 (
            .O(N__15975),
            .I(N__15955));
    InMux I__2599 (
            .O(N__15974),
            .I(N__15955));
    InMux I__2598 (
            .O(N__15973),
            .I(N__15955));
    InMux I__2597 (
            .O(N__15972),
            .I(N__15955));
    LocalMux I__2596 (
            .O(N__15955),
            .I(N__15951));
    InMux I__2595 (
            .O(N__15954),
            .I(N__15948));
    Odrv4 I__2594 (
            .O(N__15951),
            .I(\buart.Z_rx.N_27_0_i ));
    LocalMux I__2593 (
            .O(N__15948),
            .I(\buart.Z_rx.N_27_0_i ));
    CascadeMux I__2592 (
            .O(N__15943),
            .I(N__15938));
    CascadeMux I__2591 (
            .O(N__15942),
            .I(N__15935));
    CascadeMux I__2590 (
            .O(N__15941),
            .I(N__15932));
    InMux I__2589 (
            .O(N__15938),
            .I(N__15902));
    InMux I__2588 (
            .O(N__15935),
            .I(N__15902));
    InMux I__2587 (
            .O(N__15932),
            .I(N__15902));
    InMux I__2586 (
            .O(N__15931),
            .I(N__15902));
    InMux I__2585 (
            .O(N__15930),
            .I(N__15902));
    InMux I__2584 (
            .O(N__15929),
            .I(N__15902));
    InMux I__2583 (
            .O(N__15928),
            .I(N__15902));
    InMux I__2582 (
            .O(N__15927),
            .I(N__15902));
    InMux I__2581 (
            .O(N__15926),
            .I(N__15897));
    InMux I__2580 (
            .O(N__15925),
            .I(N__15897));
    InMux I__2579 (
            .O(N__15924),
            .I(N__15892));
    InMux I__2578 (
            .O(N__15923),
            .I(N__15892));
    InMux I__2577 (
            .O(N__15922),
            .I(N__15887));
    InMux I__2576 (
            .O(N__15921),
            .I(N__15887));
    InMux I__2575 (
            .O(N__15920),
            .I(N__15882));
    InMux I__2574 (
            .O(N__15919),
            .I(N__15882));
    LocalMux I__2573 (
            .O(N__15902),
            .I(\buart.Z_rx.startbit ));
    LocalMux I__2572 (
            .O(N__15897),
            .I(\buart.Z_rx.startbit ));
    LocalMux I__2571 (
            .O(N__15892),
            .I(\buart.Z_rx.startbit ));
    LocalMux I__2570 (
            .O(N__15887),
            .I(\buart.Z_rx.startbit ));
    LocalMux I__2569 (
            .O(N__15882),
            .I(\buart.Z_rx.startbit ));
    CEMux I__2568 (
            .O(N__15871),
            .I(N__15867));
    CEMux I__2567 (
            .O(N__15870),
            .I(N__15864));
    LocalMux I__2566 (
            .O(N__15867),
            .I(N__15861));
    LocalMux I__2565 (
            .O(N__15864),
            .I(N__15858));
    Span4Mux_h I__2564 (
            .O(N__15861),
            .I(N__15855));
    Span4Mux_h I__2563 (
            .O(N__15858),
            .I(N__15852));
    Span4Mux_s1_v I__2562 (
            .O(N__15855),
            .I(N__15849));
    Odrv4 I__2561 (
            .O(N__15852),
            .I(\buart.Z_rx.bitcounte_0_0 ));
    Odrv4 I__2560 (
            .O(N__15849),
            .I(\buart.Z_rx.bitcounte_0_0 ));
    InMux I__2559 (
            .O(N__15844),
            .I(N__15839));
    CascadeMux I__2558 (
            .O(N__15843),
            .I(N__15832));
    InMux I__2557 (
            .O(N__15842),
            .I(N__15829));
    LocalMux I__2556 (
            .O(N__15839),
            .I(N__15826));
    InMux I__2555 (
            .O(N__15838),
            .I(N__15817));
    InMux I__2554 (
            .O(N__15837),
            .I(N__15817));
    InMux I__2553 (
            .O(N__15836),
            .I(N__15817));
    InMux I__2552 (
            .O(N__15835),
            .I(N__15817));
    InMux I__2551 (
            .O(N__15832),
            .I(N__15814));
    LocalMux I__2550 (
            .O(N__15829),
            .I(buart__rx_bitcount_0));
    Odrv4 I__2549 (
            .O(N__15826),
            .I(buart__rx_bitcount_0));
    LocalMux I__2548 (
            .O(N__15817),
            .I(buart__rx_bitcount_0));
    LocalMux I__2547 (
            .O(N__15814),
            .I(buart__rx_bitcount_0));
    InMux I__2546 (
            .O(N__15805),
            .I(N__15800));
    CascadeMux I__2545 (
            .O(N__15804),
            .I(N__15797));
    InMux I__2544 (
            .O(N__15803),
            .I(N__15790));
    LocalMux I__2543 (
            .O(N__15800),
            .I(N__15787));
    InMux I__2542 (
            .O(N__15797),
            .I(N__15784));
    InMux I__2541 (
            .O(N__15796),
            .I(N__15781));
    InMux I__2540 (
            .O(N__15795),
            .I(N__15778));
    InMux I__2539 (
            .O(N__15794),
            .I(N__15773));
    InMux I__2538 (
            .O(N__15793),
            .I(N__15773));
    LocalMux I__2537 (
            .O(N__15790),
            .I(buart__rx_bitcount_1));
    Odrv4 I__2536 (
            .O(N__15787),
            .I(buart__rx_bitcount_1));
    LocalMux I__2535 (
            .O(N__15784),
            .I(buart__rx_bitcount_1));
    LocalMux I__2534 (
            .O(N__15781),
            .I(buart__rx_bitcount_1));
    LocalMux I__2533 (
            .O(N__15778),
            .I(buart__rx_bitcount_1));
    LocalMux I__2532 (
            .O(N__15773),
            .I(buart__rx_bitcount_1));
    CascadeMux I__2531 (
            .O(N__15760),
            .I(N__15757));
    InMux I__2530 (
            .O(N__15757),
            .I(N__15754));
    LocalMux I__2529 (
            .O(N__15754),
            .I(N__15751));
    Odrv4 I__2528 (
            .O(N__15751),
            .I(\buart.Z_rx.bitcount_cry_0_THRU_CO ));
    InMux I__2527 (
            .O(N__15748),
            .I(\buart.Z_rx.bitcount_cry_0 ));
    CascadeMux I__2526 (
            .O(N__15745),
            .I(N__15741));
    CascadeMux I__2525 (
            .O(N__15744),
            .I(N__15737));
    InMux I__2524 (
            .O(N__15741),
            .I(N__15730));
    InMux I__2523 (
            .O(N__15740),
            .I(N__15730));
    InMux I__2522 (
            .O(N__15737),
            .I(N__15730));
    LocalMux I__2521 (
            .O(N__15730),
            .I(N__15727));
    Odrv4 I__2520 (
            .O(N__15727),
            .I(\buart.Z_rx.bitcount_cry_1_THRU_CO ));
    InMux I__2519 (
            .O(N__15724),
            .I(\buart.Z_rx.bitcount_cry_1 ));
    CascadeMux I__2518 (
            .O(N__15721),
            .I(N__15717));
    InMux I__2517 (
            .O(N__15720),
            .I(N__15712));
    InMux I__2516 (
            .O(N__15717),
            .I(N__15712));
    LocalMux I__2515 (
            .O(N__15712),
            .I(N__15709));
    Odrv4 I__2514 (
            .O(N__15709),
            .I(\buart.Z_rx.bitcount_cry_2_THRU_CO ));
    InMux I__2513 (
            .O(N__15706),
            .I(\buart.Z_rx.bitcount_cry_2 ));
    InMux I__2512 (
            .O(N__15703),
            .I(\buart.Z_rx.bitcount_cry_3 ));
    CascadeMux I__2511 (
            .O(N__15700),
            .I(N__15696));
    InMux I__2510 (
            .O(N__15699),
            .I(N__15691));
    InMux I__2509 (
            .O(N__15696),
            .I(N__15691));
    LocalMux I__2508 (
            .O(N__15691),
            .I(N__15688));
    Odrv12 I__2507 (
            .O(N__15688),
            .I(\buart.Z_rx.bitcount_cry_3_THRU_CO ));
    CascadeMux I__2506 (
            .O(N__15685),
            .I(N__15682));
    InMux I__2505 (
            .O(N__15682),
            .I(N__15676));
    InMux I__2504 (
            .O(N__15681),
            .I(N__15676));
    LocalMux I__2503 (
            .O(N__15676),
            .I(buart__rx_bitcount_fast_4));
    InMux I__2502 (
            .O(N__15673),
            .I(N__15670));
    LocalMux I__2501 (
            .O(N__15670),
            .I(N__15666));
    InMux I__2500 (
            .O(N__15669),
            .I(N__15663));
    Odrv4 I__2499 (
            .O(N__15666),
            .I(buart__rx_bitcount_fast_3));
    LocalMux I__2498 (
            .O(N__15663),
            .I(buart__rx_bitcount_fast_3));
    InMux I__2497 (
            .O(N__15658),
            .I(N__15655));
    LocalMux I__2496 (
            .O(N__15655),
            .I(\Lab_UT.dictrl.decoder.g0_6_1 ));
    CascadeMux I__2495 (
            .O(N__15652),
            .I(\buart.Z_rx.un1_sample_0_cascade_ ));
    IoInMux I__2494 (
            .O(N__15649),
            .I(N__15646));
    LocalMux I__2493 (
            .O(N__15646),
            .I(N__15643));
    Odrv4 I__2492 (
            .O(N__15643),
            .I(\buart.Z_rx.sample ));
    CascadeMux I__2491 (
            .O(N__15640),
            .I(\buart.Z_rx.idle_0_cascade_ ));
    InMux I__2490 (
            .O(N__15637),
            .I(N__15633));
    InMux I__2489 (
            .O(N__15636),
            .I(N__15630));
    LocalMux I__2488 (
            .O(N__15633),
            .I(\buart.Z_rx.idle ));
    LocalMux I__2487 (
            .O(N__15630),
            .I(\buart.Z_rx.idle ));
    CascadeMux I__2486 (
            .O(N__15625),
            .I(N__15621));
    InMux I__2485 (
            .O(N__15624),
            .I(N__15616));
    InMux I__2484 (
            .O(N__15621),
            .I(N__15613));
    InMux I__2483 (
            .O(N__15620),
            .I(N__15608));
    InMux I__2482 (
            .O(N__15619),
            .I(N__15608));
    LocalMux I__2481 (
            .O(N__15616),
            .I(\buart.Z_rx.ser_clk ));
    LocalMux I__2480 (
            .O(N__15613),
            .I(\buart.Z_rx.ser_clk ));
    LocalMux I__2479 (
            .O(N__15608),
            .I(\buart.Z_rx.ser_clk ));
    CascadeMux I__2478 (
            .O(N__15601),
            .I(\buart.Z_rx.idle_cascade_ ));
    CascadeMux I__2477 (
            .O(N__15598),
            .I(Lab_UT_dictrl_decoder_de_cr_1_cascade_));
    InMux I__2476 (
            .O(N__15595),
            .I(N__15592));
    LocalMux I__2475 (
            .O(N__15592),
            .I(\Lab_UT.dictrl.N_30 ));
    InMux I__2474 (
            .O(N__15589),
            .I(N__15586));
    LocalMux I__2473 (
            .O(N__15586),
            .I(\Lab_UT.dictrl.N_41_mux ));
    CascadeMux I__2472 (
            .O(N__15583),
            .I(N__15579));
    InMux I__2471 (
            .O(N__15582),
            .I(N__15576));
    InMux I__2470 (
            .O(N__15579),
            .I(N__15572));
    LocalMux I__2469 (
            .O(N__15576),
            .I(N__15569));
    CascadeMux I__2468 (
            .O(N__15575),
            .I(N__15565));
    LocalMux I__2467 (
            .O(N__15572),
            .I(N__15562));
    Span4Mux_h I__2466 (
            .O(N__15569),
            .I(N__15559));
    InMux I__2465 (
            .O(N__15568),
            .I(N__15554));
    InMux I__2464 (
            .O(N__15565),
            .I(N__15554));
    Span4Mux_h I__2463 (
            .O(N__15562),
            .I(N__15551));
    Odrv4 I__2462 (
            .O(N__15559),
            .I(\Lab_UT.dictrl.N_34 ));
    LocalMux I__2461 (
            .O(N__15554),
            .I(\Lab_UT.dictrl.N_34 ));
    Odrv4 I__2460 (
            .O(N__15551),
            .I(\Lab_UT.dictrl.N_34 ));
    CascadeMux I__2459 (
            .O(N__15544),
            .I(\Lab_UT.dictrl.N_31_cascade_ ));
    InMux I__2458 (
            .O(N__15541),
            .I(N__15538));
    LocalMux I__2457 (
            .O(N__15538),
            .I(N__15534));
    InMux I__2456 (
            .O(N__15537),
            .I(N__15531));
    Span4Mux_s2_h I__2455 (
            .O(N__15534),
            .I(N__15528));
    LocalMux I__2454 (
            .O(N__15531),
            .I(N__15525));
    Span4Mux_v I__2453 (
            .O(N__15528),
            .I(N__15522));
    Odrv12 I__2452 (
            .O(N__15525),
            .I(\Lab_UT.dictrl.nextState_0_2 ));
    Odrv4 I__2451 (
            .O(N__15522),
            .I(\Lab_UT.dictrl.nextState_0_2 ));
    CEMux I__2450 (
            .O(N__15517),
            .I(N__15514));
    LocalMux I__2449 (
            .O(N__15514),
            .I(N__15510));
    CEMux I__2448 (
            .O(N__15513),
            .I(N__15507));
    Span4Mux_v I__2447 (
            .O(N__15510),
            .I(N__15504));
    LocalMux I__2446 (
            .O(N__15507),
            .I(N__15501));
    Odrv4 I__2445 (
            .O(N__15504),
            .I(\Lab_UT.dictrl.currState_0_ret_29_RNIDFRSEEZ0 ));
    Odrv12 I__2444 (
            .O(N__15501),
            .I(\Lab_UT.dictrl.currState_0_ret_29_RNIDFRSEEZ0 ));
    CascadeMux I__2443 (
            .O(N__15496),
            .I(N__15493));
    InMux I__2442 (
            .O(N__15493),
            .I(N__15490));
    LocalMux I__2441 (
            .O(N__15490),
            .I(buart__rx_bitcount_fast_2));
    CascadeMux I__2440 (
            .O(N__15487),
            .I(\Lab_UT.dictrl.r_dicLdMtens20_0_cascade_ ));
    InMux I__2439 (
            .O(N__15484),
            .I(N__15477));
    InMux I__2438 (
            .O(N__15483),
            .I(N__15467));
    InMux I__2437 (
            .O(N__15482),
            .I(N__15467));
    InMux I__2436 (
            .O(N__15481),
            .I(N__15462));
    InMux I__2435 (
            .O(N__15480),
            .I(N__15462));
    LocalMux I__2434 (
            .O(N__15477),
            .I(N__15459));
    InMux I__2433 (
            .O(N__15476),
            .I(N__15456));
    InMux I__2432 (
            .O(N__15475),
            .I(N__15451));
    InMux I__2431 (
            .O(N__15474),
            .I(N__15451));
    InMux I__2430 (
            .O(N__15473),
            .I(N__15446));
    InMux I__2429 (
            .O(N__15472),
            .I(N__15446));
    LocalMux I__2428 (
            .O(N__15467),
            .I(N__15443));
    LocalMux I__2427 (
            .O(N__15462),
            .I(N__15440));
    Span4Mux_h I__2426 (
            .O(N__15459),
            .I(N__15435));
    LocalMux I__2425 (
            .O(N__15456),
            .I(N__15435));
    LocalMux I__2424 (
            .O(N__15451),
            .I(N__15429));
    LocalMux I__2423 (
            .O(N__15446),
            .I(N__15429));
    Span4Mux_s3_h I__2422 (
            .O(N__15443),
            .I(N__15424));
    Span4Mux_h I__2421 (
            .O(N__15440),
            .I(N__15424));
    Span4Mux_h I__2420 (
            .O(N__15435),
            .I(N__15421));
    InMux I__2419 (
            .O(N__15434),
            .I(N__15418));
    Odrv12 I__2418 (
            .O(N__15429),
            .I(\Lab_UT.dictrl.N_6ctr ));
    Odrv4 I__2417 (
            .O(N__15424),
            .I(\Lab_UT.dictrl.N_6ctr ));
    Odrv4 I__2416 (
            .O(N__15421),
            .I(\Lab_UT.dictrl.N_6ctr ));
    LocalMux I__2415 (
            .O(N__15418),
            .I(\Lab_UT.dictrl.N_6ctr ));
    InMux I__2414 (
            .O(N__15409),
            .I(N__15406));
    LocalMux I__2413 (
            .O(N__15406),
            .I(\Lab_UT.dictrl.r_dicLdMtens22_2_reti ));
    InMux I__2412 (
            .O(N__15403),
            .I(N__15400));
    LocalMux I__2411 (
            .O(N__15400),
            .I(N__15397));
    Odrv12 I__2410 (
            .O(N__15397),
            .I(\Lab_UT.dictrl.N_7_1_0 ));
    CascadeMux I__2409 (
            .O(N__15394),
            .I(\Lab_UT.dictrl.r_dicLdMtens22_2_reti_cascade_ ));
    InMux I__2408 (
            .O(N__15391),
            .I(N__15388));
    LocalMux I__2407 (
            .O(N__15388),
            .I(\Lab_UT.dictrl.g0_0_3 ));
    InMux I__2406 (
            .O(N__15385),
            .I(N__15381));
    InMux I__2405 (
            .O(N__15384),
            .I(N__15378));
    LocalMux I__2404 (
            .O(N__15381),
            .I(N__15374));
    LocalMux I__2403 (
            .O(N__15378),
            .I(N__15371));
    InMux I__2402 (
            .O(N__15377),
            .I(N__15368));
    Span4Mux_h I__2401 (
            .O(N__15374),
            .I(N__15363));
    Span4Mux_v I__2400 (
            .O(N__15371),
            .I(N__15363));
    LocalMux I__2399 (
            .O(N__15368),
            .I(\Lab_UT.dictrl.N_10ctr ));
    Odrv4 I__2398 (
            .O(N__15363),
            .I(\Lab_UT.dictrl.N_10ctr ));
    InMux I__2397 (
            .O(N__15358),
            .I(N__15352));
    InMux I__2396 (
            .O(N__15357),
            .I(N__15352));
    LocalMux I__2395 (
            .O(N__15352),
            .I(\Lab_UT.dictrl.r_dicLdMtens22_4_0 ));
    InMux I__2394 (
            .O(N__15349),
            .I(N__15346));
    LocalMux I__2393 (
            .O(N__15346),
            .I(N__15343));
    Span4Mux_h I__2392 (
            .O(N__15343),
            .I(N__15340));
    Odrv4 I__2391 (
            .O(N__15340),
            .I(N_7));
    CascadeMux I__2390 (
            .O(N__15337),
            .I(N__15333));
    InMux I__2389 (
            .O(N__15336),
            .I(N__15330));
    InMux I__2388 (
            .O(N__15333),
            .I(N__15327));
    LocalMux I__2387 (
            .O(N__15330),
            .I(N__15324));
    LocalMux I__2386 (
            .O(N__15327),
            .I(N__15321));
    Span4Mux_s3_h I__2385 (
            .O(N__15324),
            .I(N__15317));
    Span4Mux_h I__2384 (
            .O(N__15321),
            .I(N__15314));
    InMux I__2383 (
            .O(N__15320),
            .I(N__15311));
    Odrv4 I__2382 (
            .O(N__15317),
            .I(\Lab_UT.dictrl.N_20 ));
    Odrv4 I__2381 (
            .O(N__15314),
            .I(\Lab_UT.dictrl.N_20 ));
    LocalMux I__2380 (
            .O(N__15311),
            .I(\Lab_UT.dictrl.N_20 ));
    InMux I__2379 (
            .O(N__15304),
            .I(N__15301));
    LocalMux I__2378 (
            .O(N__15301),
            .I(N__15298));
    Span4Mux_h I__2377 (
            .O(N__15298),
            .I(N__15294));
    InMux I__2376 (
            .O(N__15297),
            .I(N__15291));
    Odrv4 I__2375 (
            .O(N__15294),
            .I(\Lab_UT.dictrl.de_littleA ));
    LocalMux I__2374 (
            .O(N__15291),
            .I(\Lab_UT.dictrl.de_littleA ));
    CascadeMux I__2373 (
            .O(N__15286),
            .I(\Lab_UT.dictrl.g2_cascade_ ));
    CascadeMux I__2372 (
            .O(N__15283),
            .I(\Lab_UT.dictrl.nextState_RNO_9Z0Z_1_cascade_ ));
    InMux I__2371 (
            .O(N__15280),
            .I(N__15276));
    InMux I__2370 (
            .O(N__15279),
            .I(N__15273));
    LocalMux I__2369 (
            .O(N__15276),
            .I(N__15268));
    LocalMux I__2368 (
            .O(N__15273),
            .I(N__15268));
    Span4Mux_v I__2367 (
            .O(N__15268),
            .I(N__15265));
    Odrv4 I__2366 (
            .O(N__15265),
            .I(\Lab_UT.dictrl.g0_i_a4_1 ));
    CascadeMux I__2365 (
            .O(N__15262),
            .I(\Lab_UT.dictrl.nextState_RNO_4Z0Z_1_cascade_ ));
    InMux I__2364 (
            .O(N__15259),
            .I(N__15256));
    LocalMux I__2363 (
            .O(N__15256),
            .I(\Lab_UT.dictrl.nextState_RNO_3Z0Z_1 ));
    InMux I__2362 (
            .O(N__15253),
            .I(N__15250));
    LocalMux I__2361 (
            .O(N__15250),
            .I(N__15247));
    Odrv12 I__2360 (
            .O(N__15247),
            .I(\Lab_UT.dictrl.g0_i_o4_5 ));
    InMux I__2359 (
            .O(N__15244),
            .I(N__15241));
    LocalMux I__2358 (
            .O(N__15241),
            .I(\Lab_UT.dictrl.N_11 ));
    InMux I__2357 (
            .O(N__15238),
            .I(N__15235));
    LocalMux I__2356 (
            .O(N__15235),
            .I(\Lab_UT.dictrl.N_18_0 ));
    CascadeMux I__2355 (
            .O(N__15232),
            .I(N__15229));
    InMux I__2354 (
            .O(N__15229),
            .I(N__15226));
    LocalMux I__2353 (
            .O(N__15226),
            .I(\Lab_UT.dictrl.g1_3_0 ));
    InMux I__2352 (
            .O(N__15223),
            .I(N__15220));
    LocalMux I__2351 (
            .O(N__15220),
            .I(N__15217));
    Odrv4 I__2350 (
            .O(N__15217),
            .I(\Lab_UT.dictrl.N_13_0 ));
    CascadeMux I__2349 (
            .O(N__15214),
            .I(\Lab_UT.dictrl.g1_4_0_cascade_ ));
    InMux I__2348 (
            .O(N__15211),
            .I(N__15208));
    LocalMux I__2347 (
            .O(N__15208),
            .I(\Lab_UT.dictrl.N_14 ));
    CascadeMux I__2346 (
            .O(N__15205),
            .I(\Lab_UT.dictrl.N_36_0_cascade_ ));
    CascadeMux I__2345 (
            .O(N__15202),
            .I(\Lab_UT.dictrl.nextStateZ0Z_3_cascade_ ));
    InMux I__2344 (
            .O(N__15199),
            .I(N__15196));
    LocalMux I__2343 (
            .O(N__15196),
            .I(\Lab_UT.dictrl.r_dicLdMtens21_1 ));
    InMux I__2342 (
            .O(N__15193),
            .I(N__15189));
    InMux I__2341 (
            .O(N__15192),
            .I(N__15186));
    LocalMux I__2340 (
            .O(N__15189),
            .I(\Lab_UT.dictrl.N_18 ));
    LocalMux I__2339 (
            .O(N__15186),
            .I(\Lab_UT.dictrl.N_18 ));
    InMux I__2338 (
            .O(N__15181),
            .I(N__15178));
    LocalMux I__2337 (
            .O(N__15178),
            .I(\Lab_UT.dictrl.N_33 ));
    InMux I__2336 (
            .O(N__15175),
            .I(N__15172));
    LocalMux I__2335 (
            .O(N__15172),
            .I(\Lab_UT.dictrl.N_1607_0_0 ));
    InMux I__2334 (
            .O(N__15169),
            .I(N__15166));
    LocalMux I__2333 (
            .O(N__15166),
            .I(\Lab_UT.dictrl.N_10_0_0 ));
    InMux I__2332 (
            .O(N__15163),
            .I(N__15160));
    LocalMux I__2331 (
            .O(N__15160),
            .I(\Lab_UT.dictrl.g1 ));
    CascadeMux I__2330 (
            .O(N__15157),
            .I(N__15154));
    InMux I__2329 (
            .O(N__15154),
            .I(N__15151));
    LocalMux I__2328 (
            .O(N__15151),
            .I(N__15148));
    Span4Mux_h I__2327 (
            .O(N__15148),
            .I(N__15145));
    Odrv4 I__2326 (
            .O(N__15145),
            .I(\Lab_UT.dictrl.N_1614_0 ));
    CascadeMux I__2325 (
            .O(N__15142),
            .I(N__15139));
    InMux I__2324 (
            .O(N__15139),
            .I(N__15136));
    LocalMux I__2323 (
            .O(N__15136),
            .I(\Lab_UT.dictrl.N_26 ));
    InMux I__2322 (
            .O(N__15133),
            .I(N__15130));
    LocalMux I__2321 (
            .O(N__15130),
            .I(\Lab_UT.dictrl.un1_currState_6 ));
    InMux I__2320 (
            .O(N__15127),
            .I(N__15121));
    InMux I__2319 (
            .O(N__15126),
            .I(N__15121));
    LocalMux I__2318 (
            .O(N__15121),
            .I(\Lab_UT.dictrl.r_enableZ0Z1 ));
    InMux I__2317 (
            .O(N__15118),
            .I(N__15112));
    InMux I__2316 (
            .O(N__15117),
            .I(N__15112));
    LocalMux I__2315 (
            .O(N__15112),
            .I(N__15104));
    InMux I__2314 (
            .O(N__15111),
            .I(N__15099));
    InMux I__2313 (
            .O(N__15110),
            .I(N__15099));
    InMux I__2312 (
            .O(N__15109),
            .I(N__15096));
    InMux I__2311 (
            .O(N__15108),
            .I(N__15091));
    InMux I__2310 (
            .O(N__15107),
            .I(N__15091));
    Sp12to4 I__2309 (
            .O(N__15104),
            .I(N__15088));
    LocalMux I__2308 (
            .O(N__15099),
            .I(N__15081));
    LocalMux I__2307 (
            .O(N__15096),
            .I(N__15081));
    LocalMux I__2306 (
            .O(N__15091),
            .I(N__15081));
    Odrv12 I__2305 (
            .O(N__15088),
            .I(\Lab_UT.dictrl.enableSeg3 ));
    Odrv4 I__2304 (
            .O(N__15081),
            .I(\Lab_UT.dictrl.enableSeg3 ));
    CascadeMux I__2303 (
            .O(N__15076),
            .I(N__15073));
    InMux I__2302 (
            .O(N__15073),
            .I(N__15067));
    InMux I__2301 (
            .O(N__15072),
            .I(N__15067));
    LocalMux I__2300 (
            .O(N__15067),
            .I(\Lab_UT.dictrl.r_enableZ0Z3 ));
    CascadeMux I__2299 (
            .O(N__15064),
            .I(N__15061));
    InMux I__2298 (
            .O(N__15061),
            .I(N__15056));
    InMux I__2297 (
            .O(N__15060),
            .I(N__15050));
    InMux I__2296 (
            .O(N__15059),
            .I(N__15050));
    LocalMux I__2295 (
            .O(N__15056),
            .I(N__15047));
    InMux I__2294 (
            .O(N__15055),
            .I(N__15044));
    LocalMux I__2293 (
            .O(N__15050),
            .I(N__15041));
    Span4Mux_v I__2292 (
            .O(N__15047),
            .I(N__15035));
    LocalMux I__2291 (
            .O(N__15044),
            .I(N__15032));
    Span4Mux_h I__2290 (
            .O(N__15041),
            .I(N__15029));
    InMux I__2289 (
            .O(N__15040),
            .I(N__15022));
    InMux I__2288 (
            .O(N__15039),
            .I(N__15022));
    InMux I__2287 (
            .O(N__15038),
            .I(N__15022));
    Odrv4 I__2286 (
            .O(N__15035),
            .I(\Lab_UT.dictrl.enableSeg4 ));
    Odrv4 I__2285 (
            .O(N__15032),
            .I(\Lab_UT.dictrl.enableSeg4 ));
    Odrv4 I__2284 (
            .O(N__15029),
            .I(\Lab_UT.dictrl.enableSeg4 ));
    LocalMux I__2283 (
            .O(N__15022),
            .I(\Lab_UT.dictrl.enableSeg4 ));
    InMux I__2282 (
            .O(N__15013),
            .I(N__15010));
    LocalMux I__2281 (
            .O(N__15010),
            .I(N__15007));
    Odrv4 I__2280 (
            .O(N__15007),
            .I(\Lab_UT.dictrl.un1_currState_7 ));
    CascadeMux I__2279 (
            .O(N__15004),
            .I(N__15001));
    InMux I__2278 (
            .O(N__15001),
            .I(N__14995));
    InMux I__2277 (
            .O(N__15000),
            .I(N__14995));
    LocalMux I__2276 (
            .O(N__14995),
            .I(\Lab_UT.dictrl.r_enableZ0Z4 ));
    InMux I__2275 (
            .O(N__14992),
            .I(N__14989));
    LocalMux I__2274 (
            .O(N__14989),
            .I(N__14986));
    Odrv4 I__2273 (
            .O(N__14986),
            .I(\Lab_UT.dictrl.N_1605_1_0 ));
    CascadeMux I__2272 (
            .O(N__14983),
            .I(\Lab_UT.N_76_cascade_ ));
    CascadeMux I__2271 (
            .O(N__14980),
            .I(N__14977));
    InMux I__2270 (
            .O(N__14977),
            .I(N__14974));
    LocalMux I__2269 (
            .O(N__14974),
            .I(N__14971));
    Odrv4 I__2268 (
            .O(N__14971),
            .I(\uu2.bitmapZ0Z_194 ));
    CascadeMux I__2267 (
            .O(N__14968),
            .I(\Lab_UT.L3_segment4_1_1_cascade_ ));
    InMux I__2266 (
            .O(N__14965),
            .I(N__14962));
    LocalMux I__2265 (
            .O(N__14962),
            .I(N__14959));
    Odrv4 I__2264 (
            .O(N__14959),
            .I(\uu2.bitmapZ0Z_69 ));
    InMux I__2263 (
            .O(N__14956),
            .I(N__14953));
    LocalMux I__2262 (
            .O(N__14953),
            .I(\Lab_UT.L3_segment4_1_0 ));
    InMux I__2261 (
            .O(N__14950),
            .I(N__14947));
    LocalMux I__2260 (
            .O(N__14947),
            .I(N__14944));
    Odrv4 I__2259 (
            .O(N__14944),
            .I(\uu2.bitmapZ0Z_34 ));
    CascadeMux I__2258 (
            .O(N__14941),
            .I(\Lab_UT.segment_1_6_cascade_ ));
    InMux I__2257 (
            .O(N__14938),
            .I(N__14935));
    LocalMux I__2256 (
            .O(N__14935),
            .I(N__14932));
    Odrv12 I__2255 (
            .O(N__14932),
            .I(\uu2.bitmapZ0Z_162 ));
    InMux I__2254 (
            .O(N__14929),
            .I(N__14926));
    LocalMux I__2253 (
            .O(N__14926),
            .I(N__14923));
    Odrv4 I__2252 (
            .O(N__14923),
            .I(\uu2.bitmap_pmux_sn_N_15 ));
    InMux I__2251 (
            .O(N__14920),
            .I(N__14910));
    InMux I__2250 (
            .O(N__14919),
            .I(N__14910));
    InMux I__2249 (
            .O(N__14918),
            .I(N__14910));
    InMux I__2248 (
            .O(N__14917),
            .I(N__14903));
    LocalMux I__2247 (
            .O(N__14910),
            .I(N__14900));
    InMux I__2246 (
            .O(N__14909),
            .I(N__14891));
    InMux I__2245 (
            .O(N__14908),
            .I(N__14891));
    InMux I__2244 (
            .O(N__14907),
            .I(N__14891));
    InMux I__2243 (
            .O(N__14906),
            .I(N__14888));
    LocalMux I__2242 (
            .O(N__14903),
            .I(N__14885));
    Span4Mux_h I__2241 (
            .O(N__14900),
            .I(N__14882));
    InMux I__2240 (
            .O(N__14899),
            .I(N__14877));
    InMux I__2239 (
            .O(N__14898),
            .I(N__14877));
    LocalMux I__2238 (
            .O(N__14891),
            .I(N__14874));
    LocalMux I__2237 (
            .O(N__14888),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    Odrv12 I__2236 (
            .O(N__14885),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    Odrv4 I__2235 (
            .O(N__14882),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    LocalMux I__2234 (
            .O(N__14877),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    Odrv4 I__2233 (
            .O(N__14874),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    InMux I__2232 (
            .O(N__14863),
            .I(N__14860));
    LocalMux I__2231 (
            .O(N__14860),
            .I(N__14857));
    Odrv4 I__2230 (
            .O(N__14857),
            .I(\Lab_UT.L3_segment3_0_i_1_0 ));
    InMux I__2229 (
            .O(N__14854),
            .I(N__14851));
    LocalMux I__2228 (
            .O(N__14851),
            .I(N__14848));
    Odrv4 I__2227 (
            .O(N__14848),
            .I(\Lab_UT.L3_segment3_0_i_1_3 ));
    CascadeMux I__2226 (
            .O(N__14845),
            .I(\Lab_UT.L3_segment3_1_2_cascade_ ));
    InMux I__2225 (
            .O(N__14842),
            .I(N__14826));
    InMux I__2224 (
            .O(N__14841),
            .I(N__14826));
    InMux I__2223 (
            .O(N__14840),
            .I(N__14826));
    InMux I__2222 (
            .O(N__14839),
            .I(N__14826));
    InMux I__2221 (
            .O(N__14838),
            .I(N__14817));
    InMux I__2220 (
            .O(N__14837),
            .I(N__14817));
    InMux I__2219 (
            .O(N__14836),
            .I(N__14817));
    InMux I__2218 (
            .O(N__14835),
            .I(N__14817));
    LocalMux I__2217 (
            .O(N__14826),
            .I(\Lab_UT.Mone_at_0 ));
    LocalMux I__2216 (
            .O(N__14817),
            .I(\Lab_UT.Mone_at_0 ));
    CascadeMux I__2215 (
            .O(N__14812),
            .I(N__14805));
    CascadeMux I__2214 (
            .O(N__14811),
            .I(N__14800));
    CascadeMux I__2213 (
            .O(N__14810),
            .I(N__14797));
    InMux I__2212 (
            .O(N__14809),
            .I(N__14786));
    InMux I__2211 (
            .O(N__14808),
            .I(N__14786));
    InMux I__2210 (
            .O(N__14805),
            .I(N__14786));
    InMux I__2209 (
            .O(N__14804),
            .I(N__14786));
    InMux I__2208 (
            .O(N__14803),
            .I(N__14777));
    InMux I__2207 (
            .O(N__14800),
            .I(N__14777));
    InMux I__2206 (
            .O(N__14797),
            .I(N__14777));
    InMux I__2205 (
            .O(N__14796),
            .I(N__14777));
    InMux I__2204 (
            .O(N__14795),
            .I(N__14774));
    LocalMux I__2203 (
            .O(N__14786),
            .I(\Lab_UT.Mone_at_3 ));
    LocalMux I__2202 (
            .O(N__14777),
            .I(\Lab_UT.Mone_at_3 ));
    LocalMux I__2201 (
            .O(N__14774),
            .I(\Lab_UT.Mone_at_3 ));
    CascadeMux I__2200 (
            .O(N__14767),
            .I(N__14758));
    CascadeMux I__2199 (
            .O(N__14766),
            .I(N__14755));
    CascadeMux I__2198 (
            .O(N__14765),
            .I(N__14751));
    InMux I__2197 (
            .O(N__14764),
            .I(N__14742));
    InMux I__2196 (
            .O(N__14763),
            .I(N__14742));
    InMux I__2195 (
            .O(N__14762),
            .I(N__14742));
    InMux I__2194 (
            .O(N__14761),
            .I(N__14742));
    InMux I__2193 (
            .O(N__14758),
            .I(N__14733));
    InMux I__2192 (
            .O(N__14755),
            .I(N__14733));
    InMux I__2191 (
            .O(N__14754),
            .I(N__14733));
    InMux I__2190 (
            .O(N__14751),
            .I(N__14733));
    LocalMux I__2189 (
            .O(N__14742),
            .I(\Lab_UT.Mone_at_2 ));
    LocalMux I__2188 (
            .O(N__14733),
            .I(\Lab_UT.Mone_at_2 ));
    CascadeMux I__2187 (
            .O(N__14728),
            .I(N__14724));
    CascadeMux I__2186 (
            .O(N__14727),
            .I(N__14721));
    InMux I__2185 (
            .O(N__14724),
            .I(N__14706));
    InMux I__2184 (
            .O(N__14721),
            .I(N__14706));
    InMux I__2183 (
            .O(N__14720),
            .I(N__14706));
    InMux I__2182 (
            .O(N__14719),
            .I(N__14706));
    InMux I__2181 (
            .O(N__14718),
            .I(N__14697));
    InMux I__2180 (
            .O(N__14717),
            .I(N__14697));
    InMux I__2179 (
            .O(N__14716),
            .I(N__14697));
    InMux I__2178 (
            .O(N__14715),
            .I(N__14697));
    LocalMux I__2177 (
            .O(N__14706),
            .I(\Lab_UT.Mone_at_1 ));
    LocalMux I__2176 (
            .O(N__14697),
            .I(\Lab_UT.Mone_at_1 ));
    CascadeMux I__2175 (
            .O(N__14692),
            .I(\Lab_UT.L3_segment3_1_1_cascade_ ));
    InMux I__2174 (
            .O(N__14689),
            .I(N__14686));
    LocalMux I__2173 (
            .O(N__14686),
            .I(\uu2.bitmapZ0Z_203 ));
    InMux I__2172 (
            .O(N__14683),
            .I(N__14680));
    LocalMux I__2171 (
            .O(N__14680),
            .I(\uu2.bitmapZ0Z_75 ));
    InMux I__2170 (
            .O(N__14677),
            .I(N__14674));
    LocalMux I__2169 (
            .O(N__14674),
            .I(\uu2.bitmap_pmux_24_bm_1 ));
    InMux I__2168 (
            .O(N__14671),
            .I(N__14668));
    LocalMux I__2167 (
            .O(N__14668),
            .I(N__14665));
    Span4Mux_v I__2166 (
            .O(N__14665),
            .I(N__14662));
    Odrv4 I__2165 (
            .O(N__14662),
            .I(\uu2.N_48 ));
    InMux I__2164 (
            .O(N__14659),
            .I(N__14656));
    LocalMux I__2163 (
            .O(N__14656),
            .I(\uu2.bitmap_pmux_24_am_1 ));
    InMux I__2162 (
            .O(N__14653),
            .I(N__14650));
    LocalMux I__2161 (
            .O(N__14650),
            .I(\uu2.bitmapZ0Z_87 ));
    CascadeMux I__2160 (
            .O(N__14647),
            .I(\uu2.N_386_cascade_ ));
    CascadeMux I__2159 (
            .O(N__14644),
            .I(\uu2.w_addr_displaying_nesr_RNI1JET2Z0Z_7_cascade_ ));
    InMux I__2158 (
            .O(N__14641),
            .I(N__14635));
    InMux I__2157 (
            .O(N__14640),
            .I(N__14635));
    LocalMux I__2156 (
            .O(N__14635),
            .I(\uu2.bitmapZ0Z_314 ));
    InMux I__2155 (
            .O(N__14632),
            .I(N__14629));
    LocalMux I__2154 (
            .O(N__14629),
            .I(\uu2.bitmap_pmux_23_ns_1 ));
    InMux I__2153 (
            .O(N__14626),
            .I(N__14623));
    LocalMux I__2152 (
            .O(N__14623),
            .I(\uu2.bitmap_pmux_sn_N_20 ));
    InMux I__2151 (
            .O(N__14620),
            .I(N__14617));
    LocalMux I__2150 (
            .O(N__14617),
            .I(N__14614));
    Odrv4 I__2149 (
            .O(N__14614),
            .I(\uu2.bitmapZ0Z_168 ));
    CascadeMux I__2148 (
            .O(N__14611),
            .I(\uu2.N_17_cascade_ ));
    InMux I__2147 (
            .O(N__14608),
            .I(N__14605));
    LocalMux I__2146 (
            .O(N__14605),
            .I(\uu2.bitmap_RNIELSJ2Z0Z_111 ));
    InMux I__2145 (
            .O(N__14602),
            .I(N__14599));
    LocalMux I__2144 (
            .O(N__14599),
            .I(\uu2.bitmap_pmux_sn_N_54_mux ));
    InMux I__2143 (
            .O(N__14596),
            .I(N__14593));
    LocalMux I__2142 (
            .O(N__14593),
            .I(\uu2.bitmapZ0Z_111 ));
    CascadeMux I__2141 (
            .O(N__14590),
            .I(N__14586));
    InMux I__2140 (
            .O(N__14589),
            .I(N__14578));
    InMux I__2139 (
            .O(N__14586),
            .I(N__14578));
    InMux I__2138 (
            .O(N__14585),
            .I(N__14578));
    LocalMux I__2137 (
            .O(N__14578),
            .I(N__14575));
    Span4Mux_v I__2136 (
            .O(N__14575),
            .I(N__14572));
    Odrv4 I__2135 (
            .O(N__14572),
            .I(\uu2.bitmap_pmux_sn_N_33 ));
    CascadeMux I__2134 (
            .O(N__14569),
            .I(\uu2.N_39_cascade_ ));
    CascadeMux I__2133 (
            .O(N__14566),
            .I(\resetGen.reset_count_2_0_4_cascade_ ));
    CascadeMux I__2132 (
            .O(N__14563),
            .I(N__14560));
    InMux I__2131 (
            .O(N__14560),
            .I(N__14557));
    LocalMux I__2130 (
            .O(N__14557),
            .I(N__14554));
    Odrv4 I__2129 (
            .O(N__14554),
            .I(\uu2.mem0.w_addr_2 ));
    CascadeMux I__2128 (
            .O(N__14551),
            .I(N__14548));
    InMux I__2127 (
            .O(N__14548),
            .I(N__14545));
    LocalMux I__2126 (
            .O(N__14545),
            .I(N__14542));
    Span4Mux_s3_h I__2125 (
            .O(N__14542),
            .I(N__14539));
    Odrv4 I__2124 (
            .O(N__14539),
            .I(\uu2.mem0.w_addr_4 ));
    CascadeMux I__2123 (
            .O(N__14536),
            .I(N__14533));
    InMux I__2122 (
            .O(N__14533),
            .I(N__14530));
    LocalMux I__2121 (
            .O(N__14530),
            .I(N__14527));
    Odrv4 I__2120 (
            .O(N__14527),
            .I(\uu2.mem0.w_addr_5 ));
    CascadeMux I__2119 (
            .O(N__14524),
            .I(N__14521));
    InMux I__2118 (
            .O(N__14521),
            .I(N__14518));
    LocalMux I__2117 (
            .O(N__14518),
            .I(N__14515));
    Odrv12 I__2116 (
            .O(N__14515),
            .I(\uu2.mem0.w_addr_6 ));
    CascadeMux I__2115 (
            .O(N__14512),
            .I(\Lab_UT.dictrl.decoder.g0Z0Z_7_cascade_ ));
    InMux I__2114 (
            .O(N__14509),
            .I(N__14505));
    CascadeMux I__2113 (
            .O(N__14508),
            .I(N__14502));
    LocalMux I__2112 (
            .O(N__14505),
            .I(N__14497));
    InMux I__2111 (
            .O(N__14502),
            .I(N__14494));
    InMux I__2110 (
            .O(N__14501),
            .I(N__14491));
    InMux I__2109 (
            .O(N__14500),
            .I(N__14488));
    Sp12to4 I__2108 (
            .O(N__14497),
            .I(N__14483));
    LocalMux I__2107 (
            .O(N__14494),
            .I(N__14483));
    LocalMux I__2106 (
            .O(N__14491),
            .I(N__14480));
    LocalMux I__2105 (
            .O(N__14488),
            .I(N__14477));
    Span12Mux_s5_v I__2104 (
            .O(N__14483),
            .I(N__14474));
    Odrv4 I__2103 (
            .O(N__14480),
            .I(\Lab_UT.dictrl.currState_fast_0 ));
    Odrv4 I__2102 (
            .O(N__14477),
            .I(\Lab_UT.dictrl.currState_fast_0 ));
    Odrv12 I__2101 (
            .O(N__14474),
            .I(\Lab_UT.dictrl.currState_fast_0 ));
    CascadeMux I__2100 (
            .O(N__14467),
            .I(\Lab_UT.dictrl.g1_4_1_0_cascade_ ));
    InMux I__2099 (
            .O(N__14464),
            .I(N__14461));
    LocalMux I__2098 (
            .O(N__14461),
            .I(\Lab_UT.dictrl.de_littleA_0 ));
    CascadeMux I__2097 (
            .O(N__14458),
            .I(\Lab_UT.dictrl.g1_4_cascade_ ));
    InMux I__2096 (
            .O(N__14455),
            .I(N__14452));
    LocalMux I__2095 (
            .O(N__14452),
            .I(N__14449));
    Span4Mux_v I__2094 (
            .O(N__14449),
            .I(N__14446));
    Odrv4 I__2093 (
            .O(N__14446),
            .I(\Lab_UT.dictrl.N_17_0_0 ));
    InMux I__2092 (
            .O(N__14443),
            .I(N__14440));
    LocalMux I__2091 (
            .O(N__14440),
            .I(\Lab_UT.dictrl.decoder.g0_5_1 ));
    CascadeMux I__2090 (
            .O(N__14437),
            .I(N__14434));
    InMux I__2089 (
            .O(N__14434),
            .I(N__14431));
    LocalMux I__2088 (
            .O(N__14431),
            .I(\Lab_UT.dictrl.m7_sx ));
    InMux I__2087 (
            .O(N__14428),
            .I(N__14424));
    InMux I__2086 (
            .O(N__14427),
            .I(N__14421));
    LocalMux I__2085 (
            .O(N__14424),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_3 ));
    LocalMux I__2084 (
            .O(N__14421),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_3 ));
    InMux I__2083 (
            .O(N__14416),
            .I(N__14410));
    InMux I__2082 (
            .O(N__14415),
            .I(N__14407));
    InMux I__2081 (
            .O(N__14414),
            .I(N__14402));
    InMux I__2080 (
            .O(N__14413),
            .I(N__14402));
    LocalMux I__2079 (
            .O(N__14410),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ));
    LocalMux I__2078 (
            .O(N__14407),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ));
    LocalMux I__2077 (
            .O(N__14402),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ));
    InMux I__2076 (
            .O(N__14395),
            .I(N__14392));
    LocalMux I__2075 (
            .O(N__14392),
            .I(\buart.Z_rx.Z_baudgen.ser_clk_3 ));
    InMux I__2074 (
            .O(N__14389),
            .I(N__14386));
    LocalMux I__2073 (
            .O(N__14386),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO ));
    CascadeMux I__2072 (
            .O(N__14383),
            .I(\buart.Z_rx.ser_clk_cascade_ ));
    CascadeMux I__2071 (
            .O(N__14380),
            .I(N__14376));
    InMux I__2070 (
            .O(N__14379),
            .I(N__14372));
    InMux I__2069 (
            .O(N__14376),
            .I(N__14367));
    InMux I__2068 (
            .O(N__14375),
            .I(N__14367));
    LocalMux I__2067 (
            .O(N__14372),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_4 ));
    LocalMux I__2066 (
            .O(N__14367),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_4 ));
    CascadeMux I__2065 (
            .O(N__14362),
            .I(N__14358));
    InMux I__2064 (
            .O(N__14361),
            .I(N__14353));
    InMux I__2063 (
            .O(N__14358),
            .I(N__14353));
    LocalMux I__2062 (
            .O(N__14353),
            .I(bu_rx_data_fast_7));
    CascadeMux I__2061 (
            .O(N__14350),
            .I(\Lab_UT.dictrl.decoder.g0_5_0_cascade_ ));
    InMux I__2060 (
            .O(N__14347),
            .I(N__14344));
    LocalMux I__2059 (
            .O(N__14344),
            .I(N__14341));
    Odrv4 I__2058 (
            .O(N__14341),
            .I(\Lab_UT.dictrl.de_cr_0_0 ));
    InMux I__2057 (
            .O(N__14338),
            .I(N__14335));
    LocalMux I__2056 (
            .O(N__14335),
            .I(N__14332));
    Odrv4 I__2055 (
            .O(N__14332),
            .I(\Lab_UT.dictrl.decoder.g0_6_0 ));
    InMux I__2054 (
            .O(N__14329),
            .I(N__14323));
    InMux I__2053 (
            .O(N__14328),
            .I(N__14323));
    LocalMux I__2052 (
            .O(N__14323),
            .I(bu_rx_data_fast_6));
    InMux I__2051 (
            .O(N__14320),
            .I(N__14317));
    LocalMux I__2050 (
            .O(N__14317),
            .I(\Lab_UT.dictrl.decoder.g0Z0Z_4 ));
    InMux I__2049 (
            .O(N__14314),
            .I(N__14308));
    InMux I__2048 (
            .O(N__14313),
            .I(N__14308));
    LocalMux I__2047 (
            .O(N__14308),
            .I(bu_rx_data_fast_4));
    InMux I__2046 (
            .O(N__14305),
            .I(N__14299));
    InMux I__2045 (
            .O(N__14304),
            .I(N__14299));
    LocalMux I__2044 (
            .O(N__14299),
            .I(bu_rx_data_fast_5));
    CascadeMux I__2043 (
            .O(N__14296),
            .I(N__14293));
    InMux I__2042 (
            .O(N__14293),
            .I(N__14289));
    InMux I__2041 (
            .O(N__14292),
            .I(N__14286));
    LocalMux I__2040 (
            .O(N__14289),
            .I(N__14283));
    LocalMux I__2039 (
            .O(N__14286),
            .I(N__14278));
    Span4Mux_h I__2038 (
            .O(N__14283),
            .I(N__14278));
    Odrv4 I__2037 (
            .O(N__14278),
            .I(\buart.Z_rx.hhZ0Z_0 ));
    CascadeMux I__2036 (
            .O(N__14275),
            .I(\buart.Z_rx.bitcount_fast_es_RNIAJ1GZ0Z_3_cascade_ ));
    CascadeMux I__2035 (
            .O(N__14272),
            .I(bu_rx_data_rdy_cascade_));
    CascadeMux I__2034 (
            .O(N__14269),
            .I(N__14265));
    InMux I__2033 (
            .O(N__14268),
            .I(N__14262));
    InMux I__2032 (
            .O(N__14265),
            .I(N__14259));
    LocalMux I__2031 (
            .O(N__14262),
            .I(N__14256));
    LocalMux I__2030 (
            .O(N__14259),
            .I(N__14253));
    Span4Mux_h I__2029 (
            .O(N__14256),
            .I(N__14250));
    Span4Mux_h I__2028 (
            .O(N__14253),
            .I(N__14247));
    Odrv4 I__2027 (
            .O(N__14250),
            .I(\Lab_UT.dictrl.N_5_0_1 ));
    Odrv4 I__2026 (
            .O(N__14247),
            .I(\Lab_UT.dictrl.N_5_0_1 ));
    CascadeMux I__2025 (
            .O(N__14242),
            .I(\Lab_UT.dictrl.g0_3_1_cascade_ ));
    InMux I__2024 (
            .O(N__14239),
            .I(N__14236));
    LocalMux I__2023 (
            .O(N__14236),
            .I(N__14233));
    Odrv4 I__2022 (
            .O(N__14233),
            .I(\Lab_UT.dictrl.g0_1_0_0 ));
    InMux I__2021 (
            .O(N__14230),
            .I(N__14227));
    LocalMux I__2020 (
            .O(N__14227),
            .I(bu_rx_data_fast_0));
    InMux I__2019 (
            .O(N__14224),
            .I(N__14219));
    InMux I__2018 (
            .O(N__14223),
            .I(N__14214));
    InMux I__2017 (
            .O(N__14222),
            .I(N__14214));
    LocalMux I__2016 (
            .O(N__14219),
            .I(\Lab_UT.dictrl.de_num_1_2 ));
    LocalMux I__2015 (
            .O(N__14214),
            .I(\Lab_UT.dictrl.de_num_1_2 ));
    InMux I__2014 (
            .O(N__14209),
            .I(N__14206));
    LocalMux I__2013 (
            .O(N__14206),
            .I(N__14202));
    InMux I__2012 (
            .O(N__14205),
            .I(N__14199));
    Odrv4 I__2011 (
            .O(N__14202),
            .I(\Lab_UT.dictrl.N_23_0_0 ));
    LocalMux I__2010 (
            .O(N__14199),
            .I(\Lab_UT.dictrl.N_23_0_0 ));
    InMux I__2009 (
            .O(N__14194),
            .I(N__14191));
    LocalMux I__2008 (
            .O(N__14191),
            .I(\Lab_UT.dictrl.N_13_0_0 ));
    CascadeMux I__2007 (
            .O(N__14188),
            .I(\Lab_UT.dictrl.N_14_0_0_0_cascade_ ));
    InMux I__2006 (
            .O(N__14185),
            .I(N__14182));
    LocalMux I__2005 (
            .O(N__14182),
            .I(\Lab_UT.dictrl.N_1609_0_0 ));
    InMux I__2004 (
            .O(N__14179),
            .I(N__14176));
    LocalMux I__2003 (
            .O(N__14176),
            .I(N__14172));
    InMux I__2002 (
            .O(N__14175),
            .I(N__14169));
    Span4Mux_v I__2001 (
            .O(N__14172),
            .I(N__14164));
    LocalMux I__2000 (
            .O(N__14169),
            .I(N__14164));
    Odrv4 I__1999 (
            .O(N__14164),
            .I(\Lab_UT.dictrl.N_8 ));
    InMux I__1998 (
            .O(N__14161),
            .I(N__14157));
    InMux I__1997 (
            .O(N__14160),
            .I(N__14153));
    LocalMux I__1996 (
            .O(N__14157),
            .I(N__14150));
    InMux I__1995 (
            .O(N__14156),
            .I(N__14147));
    LocalMux I__1994 (
            .O(N__14153),
            .I(\Lab_UT.dictrl.N_7 ));
    Odrv4 I__1993 (
            .O(N__14150),
            .I(\Lab_UT.dictrl.N_7 ));
    LocalMux I__1992 (
            .O(N__14147),
            .I(\Lab_UT.dictrl.N_7 ));
    CascadeMux I__1991 (
            .O(N__14140),
            .I(\Lab_UT.dictrl.N_9_0_cascade_ ));
    InMux I__1990 (
            .O(N__14137),
            .I(N__14134));
    LocalMux I__1989 (
            .O(N__14134),
            .I(\Lab_UT.dictrl.g0_6 ));
    InMux I__1988 (
            .O(N__14131),
            .I(N__14128));
    LocalMux I__1987 (
            .O(N__14128),
            .I(\Lab_UT.dictrl.N_6_0 ));
    InMux I__1986 (
            .O(N__14125),
            .I(N__14122));
    LocalMux I__1985 (
            .O(N__14122),
            .I(N__14119));
    Span4Mux_h I__1984 (
            .O(N__14119),
            .I(N__14116));
    Odrv4 I__1983 (
            .O(N__14116),
            .I(\Lab_UT.dictrl.N_9 ));
    InMux I__1982 (
            .O(N__14113),
            .I(N__14110));
    LocalMux I__1981 (
            .O(N__14110),
            .I(\Lab_UT.dictrl.m15_am ));
    InMux I__1980 (
            .O(N__14107),
            .I(N__14104));
    LocalMux I__1979 (
            .O(N__14104),
            .I(\Lab_UT.dictrl.N_20_1 ));
    InMux I__1978 (
            .O(N__14101),
            .I(N__14098));
    LocalMux I__1977 (
            .O(N__14098),
            .I(N__14092));
    CascadeMux I__1976 (
            .O(N__14097),
            .I(N__14089));
    CascadeMux I__1975 (
            .O(N__14096),
            .I(N__14084));
    CascadeMux I__1974 (
            .O(N__14095),
            .I(N__14080));
    Span4Mux_h I__1973 (
            .O(N__14092),
            .I(N__14077));
    InMux I__1972 (
            .O(N__14089),
            .I(N__14064));
    InMux I__1971 (
            .O(N__14088),
            .I(N__14064));
    InMux I__1970 (
            .O(N__14087),
            .I(N__14064));
    InMux I__1969 (
            .O(N__14084),
            .I(N__14064));
    InMux I__1968 (
            .O(N__14083),
            .I(N__14064));
    InMux I__1967 (
            .O(N__14080),
            .I(N__14064));
    Odrv4 I__1966 (
            .O(N__14077),
            .I(\Lab_UT.dictrl.currState_0_rep1 ));
    LocalMux I__1965 (
            .O(N__14064),
            .I(\Lab_UT.dictrl.currState_0_rep1 ));
    InMux I__1964 (
            .O(N__14059),
            .I(N__14056));
    LocalMux I__1963 (
            .O(N__14056),
            .I(\Lab_UT.dictrl.r_dicLdMtens17_1 ));
    CascadeMux I__1962 (
            .O(N__14053),
            .I(N__14050));
    InMux I__1961 (
            .O(N__14050),
            .I(N__14047));
    LocalMux I__1960 (
            .O(N__14047),
            .I(N__14044));
    Span4Mux_v I__1959 (
            .O(N__14044),
            .I(N__14041));
    Odrv4 I__1958 (
            .O(N__14041),
            .I(\Lab_UT.dictrl.r_dicLdMtens22_2 ));
    CascadeMux I__1957 (
            .O(N__14038),
            .I(\Lab_UT.dictrl.N_34_cascade_ ));
    InMux I__1956 (
            .O(N__14035),
            .I(N__14026));
    InMux I__1955 (
            .O(N__14034),
            .I(N__14026));
    InMux I__1954 (
            .O(N__14033),
            .I(N__14026));
    LocalMux I__1953 (
            .O(N__14026),
            .I(N__14022));
    InMux I__1952 (
            .O(N__14025),
            .I(N__14019));
    Span4Mux_h I__1951 (
            .O(N__14022),
            .I(N__14016));
    LocalMux I__1950 (
            .O(N__14019),
            .I(\Lab_UT.dictrl.currState_2_RNI0P25DZ0Z_1 ));
    Odrv4 I__1949 (
            .O(N__14016),
            .I(\Lab_UT.dictrl.currState_2_RNI0P25DZ0Z_1 ));
    CascadeMux I__1948 (
            .O(N__14011),
            .I(\Lab_UT.dictrl.m15_bm_cascade_ ));
    CascadeMux I__1947 (
            .O(N__14008),
            .I(N__14004));
    CascadeMux I__1946 (
            .O(N__14007),
            .I(N__14001));
    InMux I__1945 (
            .O(N__14004),
            .I(N__13998));
    InMux I__1944 (
            .O(N__14001),
            .I(N__13995));
    LocalMux I__1943 (
            .O(N__13998),
            .I(N__13992));
    LocalMux I__1942 (
            .O(N__13995),
            .I(\Lab_UT.dictrl.nextState_0_0 ));
    Odrv4 I__1941 (
            .O(N__13992),
            .I(\Lab_UT.dictrl.nextState_0_0 ));
    InMux I__1940 (
            .O(N__13987),
            .I(N__13984));
    LocalMux I__1939 (
            .O(N__13984),
            .I(\Lab_UT.dictrl.N_7_0 ));
    InMux I__1938 (
            .O(N__13981),
            .I(N__13978));
    LocalMux I__1937 (
            .O(N__13978),
            .I(\Lab_UT.dictrl.N_1609_1 ));
    InMux I__1936 (
            .O(N__13975),
            .I(N__13971));
    CascadeMux I__1935 (
            .O(N__13974),
            .I(N__13968));
    LocalMux I__1934 (
            .O(N__13971),
            .I(N__13965));
    InMux I__1933 (
            .O(N__13968),
            .I(N__13962));
    Odrv4 I__1932 (
            .O(N__13965),
            .I(\Lab_UT.dictrl.N_38 ));
    LocalMux I__1931 (
            .O(N__13962),
            .I(\Lab_UT.dictrl.N_38 ));
    InMux I__1930 (
            .O(N__13957),
            .I(N__13954));
    LocalMux I__1929 (
            .O(N__13954),
            .I(\Lab_UT.dictrl.currState_ret_5_RNOZ0Z_0 ));
    CascadeMux I__1928 (
            .O(N__13951),
            .I(\Lab_UT.dictrl.N_12_0_cascade_ ));
    InMux I__1927 (
            .O(N__13948),
            .I(N__13945));
    LocalMux I__1926 (
            .O(N__13945),
            .I(N__13942));
    Odrv4 I__1925 (
            .O(N__13942),
            .I(\Lab_UT.dictrl.G_28_0_a5_2_1 ));
    CascadeMux I__1924 (
            .O(N__13939),
            .I(N__13935));
    InMux I__1923 (
            .O(N__13938),
            .I(N__13932));
    InMux I__1922 (
            .O(N__13935),
            .I(N__13929));
    LocalMux I__1921 (
            .O(N__13932),
            .I(N__13926));
    LocalMux I__1920 (
            .O(N__13929),
            .I(\Lab_UT.dictrl.dicLdAMtensZ0 ));
    Odrv12 I__1919 (
            .O(N__13926),
            .I(\Lab_UT.dictrl.dicLdAMtensZ0 ));
    InMux I__1918 (
            .O(N__13921),
            .I(N__13917));
    InMux I__1917 (
            .O(N__13920),
            .I(N__13914));
    LocalMux I__1916 (
            .O(N__13917),
            .I(\Lab_UT.dictrl.dicLdAMtens_rst ));
    LocalMux I__1915 (
            .O(N__13914),
            .I(\Lab_UT.dictrl.dicLdAMtens_rst ));
    InMux I__1914 (
            .O(N__13909),
            .I(N__13906));
    LocalMux I__1913 (
            .O(N__13906),
            .I(\Lab_UT.dictrl.r_dicLdMtens16_1 ));
    CascadeMux I__1912 (
            .O(N__13903),
            .I(\Lab_UT.dictrl.g0_10_0_N_4L6_1_cascade_ ));
    SRMux I__1911 (
            .O(N__13900),
            .I(N__13897));
    LocalMux I__1910 (
            .O(N__13897),
            .I(N__13893));
    InMux I__1909 (
            .O(N__13896),
            .I(N__13890));
    Span4Mux_h I__1908 (
            .O(N__13893),
            .I(N__13887));
    LocalMux I__1907 (
            .O(N__13890),
            .I(N__13884));
    Span4Mux_v I__1906 (
            .O(N__13887),
            .I(N__13881));
    Span4Mux_h I__1905 (
            .O(N__13884),
            .I(N__13878));
    Odrv4 I__1904 (
            .O(N__13881),
            .I(\Lab_UT.dictrl.currState_ret_RNI7FNUZ0 ));
    Odrv4 I__1903 (
            .O(N__13878),
            .I(\Lab_UT.dictrl.currState_ret_RNI7FNUZ0 ));
    CascadeMux I__1902 (
            .O(N__13873),
            .I(\Lab_UT.Mone_at_0_cascade_ ));
    InMux I__1901 (
            .O(N__13870),
            .I(N__13867));
    LocalMux I__1900 (
            .O(N__13867),
            .I(\Lab_UT.N_77_0 ));
    InMux I__1899 (
            .O(N__13864),
            .I(N__13859));
    InMux I__1898 (
            .O(N__13863),
            .I(N__13854));
    InMux I__1897 (
            .O(N__13862),
            .I(N__13854));
    LocalMux I__1896 (
            .O(N__13859),
            .I(N__13851));
    LocalMux I__1895 (
            .O(N__13854),
            .I(N__13848));
    Span4Mux_h I__1894 (
            .O(N__13851),
            .I(N__13845));
    Span4Mux_h I__1893 (
            .O(N__13848),
            .I(N__13842));
    Odrv4 I__1892 (
            .O(N__13845),
            .I(\Lab_UT.dictrl.N_23 ));
    Odrv4 I__1891 (
            .O(N__13842),
            .I(\Lab_UT.dictrl.N_23 ));
    CascadeMux I__1890 (
            .O(N__13837),
            .I(\Lab_UT.dictrl.N_23_cascade_ ));
    CascadeMux I__1889 (
            .O(N__13834),
            .I(N__13831));
    InMux I__1888 (
            .O(N__13831),
            .I(N__13824));
    InMux I__1887 (
            .O(N__13830),
            .I(N__13824));
    InMux I__1886 (
            .O(N__13829),
            .I(N__13821));
    LocalMux I__1885 (
            .O(N__13824),
            .I(N__13818));
    LocalMux I__1884 (
            .O(N__13821),
            .I(N__13815));
    Span4Mux_s3_h I__1883 (
            .O(N__13818),
            .I(N__13812));
    Span4Mux_h I__1882 (
            .O(N__13815),
            .I(N__13809));
    Odrv4 I__1881 (
            .O(N__13812),
            .I(\Lab_UT.dictrl.nextState_RNIA8EV3Z0Z_1 ));
    Odrv4 I__1880 (
            .O(N__13809),
            .I(\Lab_UT.dictrl.nextState_RNIA8EV3Z0Z_1 ));
    InMux I__1879 (
            .O(N__13804),
            .I(N__13801));
    LocalMux I__1878 (
            .O(N__13801),
            .I(\Lab_UT.dictrl.N_10 ));
    CascadeMux I__1877 (
            .O(N__13798),
            .I(\Lab_UT.segmentUQ_0_0_cascade_ ));
    CascadeMux I__1876 (
            .O(N__13795),
            .I(\Lab_UT.N_65_0_cascade_ ));
    InMux I__1875 (
            .O(N__13792),
            .I(N__13789));
    LocalMux I__1874 (
            .O(N__13789),
            .I(\Lab_UT.segment_1_0_6 ));
    CascadeMux I__1873 (
            .O(N__13786),
            .I(\Lab_UT.N_76_0_cascade_ ));
    InMux I__1872 (
            .O(N__13783),
            .I(N__13780));
    LocalMux I__1871 (
            .O(N__13780),
            .I(\uu2.bitmapZ0Z_72 ));
    CascadeMux I__1870 (
            .O(N__13777),
            .I(N__13774));
    InMux I__1869 (
            .O(N__13774),
            .I(N__13771));
    LocalMux I__1868 (
            .O(N__13771),
            .I(\uu2.bitmapZ0Z_200 ));
    InMux I__1867 (
            .O(N__13768),
            .I(N__13765));
    LocalMux I__1866 (
            .O(N__13765),
            .I(\uu2.bitmap_RNIOS152Z0Z_72 ));
    InMux I__1865 (
            .O(N__13762),
            .I(N__13759));
    LocalMux I__1864 (
            .O(N__13759),
            .I(\uu2.bitmapZ0Z_40 ));
    CascadeMux I__1863 (
            .O(N__13756),
            .I(N__13753));
    InMux I__1862 (
            .O(N__13753),
            .I(N__13750));
    LocalMux I__1861 (
            .O(N__13750),
            .I(\uu2.bitmapZ0Z_296 ));
    CascadeMux I__1860 (
            .O(N__13747),
            .I(\uu2.bitmap_pmux_25_am_1_cascade_ ));
    InMux I__1859 (
            .O(N__13744),
            .I(N__13741));
    LocalMux I__1858 (
            .O(N__13741),
            .I(N__13738));
    Odrv4 I__1857 (
            .O(N__13738),
            .I(\uu2.bitmapZ0Z_197 ));
    InMux I__1856 (
            .O(N__13735),
            .I(N__13732));
    LocalMux I__1855 (
            .O(N__13732),
            .I(\uu2.bitmapZ0Z_66 ));
    CascadeMux I__1854 (
            .O(N__13729),
            .I(\uu2.bitmap_RNI2JA82Z0Z_212_cascade_ ));
    InMux I__1853 (
            .O(N__13726),
            .I(N__13722));
    InMux I__1852 (
            .O(N__13725),
            .I(N__13719));
    LocalMux I__1851 (
            .O(N__13722),
            .I(\uu2.N_31_i ));
    LocalMux I__1850 (
            .O(N__13719),
            .I(\uu2.N_31_i ));
    InMux I__1849 (
            .O(N__13714),
            .I(N__13711));
    LocalMux I__1848 (
            .O(N__13711),
            .I(\uu2.bitmap_RNIM7D32Z0Z_69 ));
    CascadeMux I__1847 (
            .O(N__13708),
            .I(\uu2.bitmap_pmux_27_ns_1_cascade_ ));
    InMux I__1846 (
            .O(N__13705),
            .I(N__13702));
    LocalMux I__1845 (
            .O(N__13702),
            .I(\uu2.N_407 ));
    CascadeMux I__1844 (
            .O(N__13699),
            .I(\uu2.un404_ci_0_cascade_ ));
    CascadeMux I__1843 (
            .O(N__13696),
            .I(N__13693));
    InMux I__1842 (
            .O(N__13693),
            .I(N__13689));
    CascadeMux I__1841 (
            .O(N__13692),
            .I(N__13685));
    LocalMux I__1840 (
            .O(N__13689),
            .I(N__13681));
    InMux I__1839 (
            .O(N__13688),
            .I(N__13674));
    InMux I__1838 (
            .O(N__13685),
            .I(N__13674));
    InMux I__1837 (
            .O(N__13684),
            .I(N__13674));
    Odrv4 I__1836 (
            .O(N__13681),
            .I(\uu2.r_addrZ0Z_6 ));
    LocalMux I__1835 (
            .O(N__13674),
            .I(\uu2.r_addrZ0Z_6 ));
    CascadeMux I__1834 (
            .O(N__13669),
            .I(N__13666));
    InMux I__1833 (
            .O(N__13666),
            .I(N__13663));
    LocalMux I__1832 (
            .O(N__13663),
            .I(N__13659));
    CascadeMux I__1831 (
            .O(N__13662),
            .I(N__13656));
    Span4Mux_h I__1830 (
            .O(N__13659),
            .I(N__13651));
    InMux I__1829 (
            .O(N__13656),
            .I(N__13648));
    InMux I__1828 (
            .O(N__13655),
            .I(N__13643));
    InMux I__1827 (
            .O(N__13654),
            .I(N__13643));
    Odrv4 I__1826 (
            .O(N__13651),
            .I(\uu2.r_addrZ0Z_2 ));
    LocalMux I__1825 (
            .O(N__13648),
            .I(\uu2.r_addrZ0Z_2 ));
    LocalMux I__1824 (
            .O(N__13643),
            .I(\uu2.r_addrZ0Z_2 ));
    CascadeMux I__1823 (
            .O(N__13636),
            .I(N__13633));
    InMux I__1822 (
            .O(N__13633),
            .I(N__13630));
    LocalMux I__1821 (
            .O(N__13630),
            .I(N__13627));
    Span4Mux_h I__1820 (
            .O(N__13627),
            .I(N__13620));
    InMux I__1819 (
            .O(N__13626),
            .I(N__13615));
    InMux I__1818 (
            .O(N__13625),
            .I(N__13615));
    InMux I__1817 (
            .O(N__13624),
            .I(N__13610));
    InMux I__1816 (
            .O(N__13623),
            .I(N__13610));
    Odrv4 I__1815 (
            .O(N__13620),
            .I(\uu2.r_addrZ0Z_1 ));
    LocalMux I__1814 (
            .O(N__13615),
            .I(\uu2.r_addrZ0Z_1 ));
    LocalMux I__1813 (
            .O(N__13610),
            .I(\uu2.r_addrZ0Z_1 ));
    CascadeMux I__1812 (
            .O(N__13603),
            .I(N__13600));
    InMux I__1811 (
            .O(N__13600),
            .I(N__13597));
    LocalMux I__1810 (
            .O(N__13597),
            .I(N__13594));
    Span4Mux_v I__1809 (
            .O(N__13594),
            .I(N__13590));
    CascadeMux I__1808 (
            .O(N__13593),
            .I(N__13586));
    Sp12to4 I__1807 (
            .O(N__13590),
            .I(N__13580));
    InMux I__1806 (
            .O(N__13589),
            .I(N__13573));
    InMux I__1805 (
            .O(N__13586),
            .I(N__13573));
    InMux I__1804 (
            .O(N__13585),
            .I(N__13573));
    InMux I__1803 (
            .O(N__13584),
            .I(N__13568));
    InMux I__1802 (
            .O(N__13583),
            .I(N__13568));
    Odrv12 I__1801 (
            .O(N__13580),
            .I(\uu2.r_addrZ0Z_0 ));
    LocalMux I__1800 (
            .O(N__13573),
            .I(\uu2.r_addrZ0Z_0 ));
    LocalMux I__1799 (
            .O(N__13568),
            .I(\uu2.r_addrZ0Z_0 ));
    CascadeMux I__1798 (
            .O(N__13561),
            .I(N__13558));
    InMux I__1797 (
            .O(N__13558),
            .I(N__13553));
    CascadeMux I__1796 (
            .O(N__13557),
            .I(N__13550));
    CascadeMux I__1795 (
            .O(N__13556),
            .I(N__13547));
    LocalMux I__1794 (
            .O(N__13553),
            .I(N__13544));
    InMux I__1793 (
            .O(N__13550),
            .I(N__13539));
    InMux I__1792 (
            .O(N__13547),
            .I(N__13539));
    Odrv4 I__1791 (
            .O(N__13544),
            .I(\uu2.r_addrZ0Z_3 ));
    LocalMux I__1790 (
            .O(N__13539),
            .I(\uu2.r_addrZ0Z_3 ));
    CEMux I__1789 (
            .O(N__13534),
            .I(N__13531));
    LocalMux I__1788 (
            .O(N__13531),
            .I(N__13528));
    Odrv12 I__1787 (
            .O(N__13528),
            .I(\uu2.trig_rd_is_det_0 ));
    CascadeMux I__1786 (
            .O(N__13525),
            .I(N__13522));
    InMux I__1785 (
            .O(N__13522),
            .I(N__13519));
    LocalMux I__1784 (
            .O(N__13519),
            .I(\uu2.bitmap_pmux_sn_N_42 ));
    CascadeMux I__1783 (
            .O(N__13516),
            .I(\uu2.bitmap_pmux_26_bm_1_cascade_ ));
    CascadeMux I__1782 (
            .O(N__13513),
            .I(N__13510));
    InMux I__1781 (
            .O(N__13510),
            .I(N__13507));
    LocalMux I__1780 (
            .O(N__13507),
            .I(\uu2.N_161 ));
    CascadeMux I__1779 (
            .O(N__13504),
            .I(\uu2.N_400_cascade_ ));
    InMux I__1778 (
            .O(N__13501),
            .I(N__13498));
    LocalMux I__1777 (
            .O(N__13498),
            .I(\uu2.N_409 ));
    InMux I__1776 (
            .O(N__13495),
            .I(N__13492));
    LocalMux I__1775 (
            .O(N__13492),
            .I(\uu2.bitmap_RNI1PH82Z0Z_34 ));
    InMux I__1774 (
            .O(N__13489),
            .I(N__13486));
    LocalMux I__1773 (
            .O(N__13486),
            .I(\uu2.N_404 ));
    InMux I__1772 (
            .O(N__13483),
            .I(N__13480));
    LocalMux I__1771 (
            .O(N__13480),
            .I(\uu2.bitmapZ0Z_290 ));
    CascadeMux I__1770 (
            .O(N__13477),
            .I(\uu2.trig_rd_is_det_cascade_ ));
    InMux I__1769 (
            .O(N__13474),
            .I(N__13471));
    LocalMux I__1768 (
            .O(N__13471),
            .I(\uu2.trig_rd_detZ0Z_1 ));
    InMux I__1767 (
            .O(N__13468),
            .I(N__13463));
    InMux I__1766 (
            .O(N__13467),
            .I(N__13460));
    InMux I__1765 (
            .O(N__13466),
            .I(N__13457));
    LocalMux I__1764 (
            .O(N__13463),
            .I(N__13454));
    LocalMux I__1763 (
            .O(N__13460),
            .I(N__13451));
    LocalMux I__1762 (
            .O(N__13457),
            .I(N__13447));
    Span4Mux_v I__1761 (
            .O(N__13454),
            .I(N__13444));
    Span4Mux_s2_v I__1760 (
            .O(N__13451),
            .I(N__13441));
    InMux I__1759 (
            .O(N__13450),
            .I(N__13438));
    Span4Mux_s3_h I__1758 (
            .O(N__13447),
            .I(N__13435));
    Odrv4 I__1757 (
            .O(N__13444),
            .I(\uu2.vram_rd_clkZ0 ));
    Odrv4 I__1756 (
            .O(N__13441),
            .I(\uu2.vram_rd_clkZ0 ));
    LocalMux I__1755 (
            .O(N__13438),
            .I(\uu2.vram_rd_clkZ0 ));
    Odrv4 I__1754 (
            .O(N__13435),
            .I(\uu2.vram_rd_clkZ0 ));
    InMux I__1753 (
            .O(N__13426),
            .I(N__13422));
    InMux I__1752 (
            .O(N__13425),
            .I(N__13419));
    LocalMux I__1751 (
            .O(N__13422),
            .I(N__13416));
    LocalMux I__1750 (
            .O(N__13419),
            .I(N__13411));
    Span4Mux_h I__1749 (
            .O(N__13416),
            .I(N__13411));
    Odrv4 I__1748 (
            .O(N__13411),
            .I(\uu2.un1_l_count_1_0 ));
    InMux I__1747 (
            .O(N__13408),
            .I(N__13402));
    InMux I__1746 (
            .O(N__13407),
            .I(N__13402));
    LocalMux I__1745 (
            .O(N__13402),
            .I(\uu2.trig_rd_detZ0Z_0 ));
    InMux I__1744 (
            .O(N__13399),
            .I(N__13396));
    LocalMux I__1743 (
            .O(N__13396),
            .I(\uu2.vbuf_raddr.un448_ci_0 ));
    CascadeMux I__1742 (
            .O(N__13393),
            .I(\uu2.vbuf_raddr.un426_ci_3_cascade_ ));
    CascadeMux I__1741 (
            .O(N__13390),
            .I(N__13387));
    InMux I__1740 (
            .O(N__13387),
            .I(N__13384));
    LocalMux I__1739 (
            .O(N__13384),
            .I(N__13380));
    InMux I__1738 (
            .O(N__13383),
            .I(N__13377));
    Span4Mux_s3_h I__1737 (
            .O(N__13380),
            .I(N__13372));
    LocalMux I__1736 (
            .O(N__13377),
            .I(N__13372));
    Odrv4 I__1735 (
            .O(N__13372),
            .I(\uu2.r_addrZ0Z_8 ));
    InMux I__1734 (
            .O(N__13369),
            .I(N__13366));
    LocalMux I__1733 (
            .O(N__13366),
            .I(\uu2.vbuf_raddr.un426_ci_3 ));
    CascadeMux I__1732 (
            .O(N__13363),
            .I(N__13360));
    InMux I__1731 (
            .O(N__13360),
            .I(N__13357));
    LocalMux I__1730 (
            .O(N__13357),
            .I(N__13352));
    InMux I__1729 (
            .O(N__13356),
            .I(N__13349));
    InMux I__1728 (
            .O(N__13355),
            .I(N__13346));
    Odrv4 I__1727 (
            .O(N__13352),
            .I(\uu2.r_addrZ0Z_7 ));
    LocalMux I__1726 (
            .O(N__13349),
            .I(\uu2.r_addrZ0Z_7 ));
    LocalMux I__1725 (
            .O(N__13346),
            .I(\uu2.r_addrZ0Z_7 ));
    InMux I__1724 (
            .O(N__13339),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_2 ));
    InMux I__1723 (
            .O(N__13336),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_3 ));
    InMux I__1722 (
            .O(N__13333),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_4 ));
    CascadeMux I__1721 (
            .O(N__13330),
            .I(N__13326));
    InMux I__1720 (
            .O(N__13329),
            .I(N__13321));
    InMux I__1719 (
            .O(N__13326),
            .I(N__13321));
    LocalMux I__1718 (
            .O(N__13321),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_5 ));
    CascadeMux I__1717 (
            .O(N__13318),
            .I(N__13315));
    InMux I__1716 (
            .O(N__13315),
            .I(N__13312));
    LocalMux I__1715 (
            .O(N__13312),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO ));
    InMux I__1714 (
            .O(N__13309),
            .I(N__13300));
    InMux I__1713 (
            .O(N__13308),
            .I(N__13300));
    InMux I__1712 (
            .O(N__13307),
            .I(N__13300));
    LocalMux I__1711 (
            .O(N__13300),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_2 ));
    CascadeMux I__1710 (
            .O(N__13297),
            .I(N__13293));
    InMux I__1709 (
            .O(N__13296),
            .I(N__13285));
    InMux I__1708 (
            .O(N__13293),
            .I(N__13285));
    InMux I__1707 (
            .O(N__13292),
            .I(N__13285));
    LocalMux I__1706 (
            .O(N__13285),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_1 ));
    CascadeMux I__1705 (
            .O(N__13282),
            .I(G_28_0_a5_0_4_cascade_));
    CascadeMux I__1704 (
            .O(N__13279),
            .I(N__13276));
    InMux I__1703 (
            .O(N__13276),
            .I(N__13273));
    LocalMux I__1702 (
            .O(N__13273),
            .I(N__13270));
    Odrv12 I__1701 (
            .O(N__13270),
            .I(shifter_RNI1D8L1_4));
    InMux I__1700 (
            .O(N__13267),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_1 ));
    CascadeMux I__1699 (
            .O(N__13264),
            .I(\Lab_UT.dictrl.decoder.g0Z0Z_5_cascade_ ));
    InMux I__1698 (
            .O(N__13261),
            .I(N__13258));
    LocalMux I__1697 (
            .O(N__13258),
            .I(\Lab_UT.dictrl.decoder.g0Z0Z_1 ));
    CascadeMux I__1696 (
            .O(N__13255),
            .I(\Lab_UT.dictrl.N_36_1_cascade_ ));
    InMux I__1695 (
            .O(N__13252),
            .I(N__13249));
    LocalMux I__1694 (
            .O(N__13249),
            .I(N__13246));
    Odrv4 I__1693 (
            .O(N__13246),
            .I(\Lab_UT.dictrl.g1_0_1 ));
    InMux I__1692 (
            .O(N__13243),
            .I(N__13240));
    LocalMux I__1691 (
            .O(N__13240),
            .I(\Lab_UT.dictrl.N_7_1 ));
    CascadeMux I__1690 (
            .O(N__13237),
            .I(N__13234));
    InMux I__1689 (
            .O(N__13234),
            .I(N__13230));
    InMux I__1688 (
            .O(N__13233),
            .I(N__13227));
    LocalMux I__1687 (
            .O(N__13230),
            .I(N__13224));
    LocalMux I__1686 (
            .O(N__13227),
            .I(N__13220));
    Span4Mux_h I__1685 (
            .O(N__13224),
            .I(N__13217));
    InMux I__1684 (
            .O(N__13223),
            .I(N__13213));
    Span4Mux_h I__1683 (
            .O(N__13220),
            .I(N__13210));
    Span4Mux_s0_h I__1682 (
            .O(N__13217),
            .I(N__13207));
    InMux I__1681 (
            .O(N__13216),
            .I(N__13204));
    LocalMux I__1680 (
            .O(N__13213),
            .I(\Lab_UT.dictrl.nextState_0_1 ));
    Odrv4 I__1679 (
            .O(N__13210),
            .I(\Lab_UT.dictrl.nextState_0_1 ));
    Odrv4 I__1678 (
            .O(N__13207),
            .I(\Lab_UT.dictrl.nextState_0_1 ));
    LocalMux I__1677 (
            .O(N__13204),
            .I(\Lab_UT.dictrl.nextState_0_1 ));
    CascadeMux I__1676 (
            .O(N__13195),
            .I(\Lab_UT.dictrl.N_20_cascade_ ));
    InMux I__1675 (
            .O(N__13192),
            .I(N__13186));
    InMux I__1674 (
            .O(N__13191),
            .I(N__13186));
    LocalMux I__1673 (
            .O(N__13186),
            .I(\Lab_UT.dictrl.G_28_0_a5_1 ));
    InMux I__1672 (
            .O(N__13183),
            .I(N__13177));
    InMux I__1671 (
            .O(N__13182),
            .I(N__13177));
    LocalMux I__1670 (
            .O(N__13177),
            .I(\Lab_UT.dictrl.N_19_0 ));
    CascadeMux I__1669 (
            .O(N__13174),
            .I(\Lab_UT.dictrl.N_8_3_cascade_ ));
    CascadeMux I__1668 (
            .O(N__13171),
            .I(\Lab_UT.dictrl.currState_2_0_rep2_RNIBGCIZ0Z9_cascade_ ));
    InMux I__1667 (
            .O(N__13168),
            .I(N__13162));
    InMux I__1666 (
            .O(N__13167),
            .I(N__13162));
    LocalMux I__1665 (
            .O(N__13162),
            .I(\Lab_UT.dictrl.G_28_0_0 ));
    InMux I__1664 (
            .O(N__13159),
            .I(N__13156));
    LocalMux I__1663 (
            .O(N__13156),
            .I(\Lab_UT.dictrl.currState_2_0_rep2_RNIKH8PZ0Z2 ));
    InMux I__1662 (
            .O(N__13153),
            .I(N__13150));
    LocalMux I__1661 (
            .O(N__13150),
            .I(shifter_RNIS6CF1_5));
    CascadeMux I__1660 (
            .O(N__13147),
            .I(\Lab_UT.dictrl.m21_rn_1_0_cascade_ ));
    InMux I__1659 (
            .O(N__13144),
            .I(N__13141));
    LocalMux I__1658 (
            .O(N__13141),
            .I(\Lab_UT.dictrl.m21_rn_0 ));
    CascadeMux I__1657 (
            .O(N__13138),
            .I(\Lab_UT.dictrl.g0_0_0_cascade_ ));
    CascadeMux I__1656 (
            .O(N__13135),
            .I(\Lab_UT.dictrl.N_1611_0_cascade_ ));
    InMux I__1655 (
            .O(N__13132),
            .I(N__13129));
    LocalMux I__1654 (
            .O(N__13129),
            .I(\Lab_UT.dictrl.N_23_0 ));
    CascadeMux I__1653 (
            .O(N__13126),
            .I(N__13123));
    InMux I__1652 (
            .O(N__13123),
            .I(N__13120));
    LocalMux I__1651 (
            .O(N__13120),
            .I(\Lab_UT.dictrl.N_8_3 ));
    InMux I__1650 (
            .O(N__13117),
            .I(N__13106));
    InMux I__1649 (
            .O(N__13116),
            .I(N__13106));
    InMux I__1648 (
            .O(N__13115),
            .I(N__13106));
    InMux I__1647 (
            .O(N__13114),
            .I(N__13103));
    InMux I__1646 (
            .O(N__13113),
            .I(N__13100));
    LocalMux I__1645 (
            .O(N__13106),
            .I(N__13097));
    LocalMux I__1644 (
            .O(N__13103),
            .I(\uu2.l_countZ0Z_1 ));
    LocalMux I__1643 (
            .O(N__13100),
            .I(\uu2.l_countZ0Z_1 ));
    Odrv4 I__1642 (
            .O(N__13097),
            .I(\uu2.l_countZ0Z_1 ));
    CascadeMux I__1641 (
            .O(N__13090),
            .I(N__13085));
    InMux I__1640 (
            .O(N__13089),
            .I(N__13080));
    InMux I__1639 (
            .O(N__13088),
            .I(N__13080));
    InMux I__1638 (
            .O(N__13085),
            .I(N__13074));
    LocalMux I__1637 (
            .O(N__13080),
            .I(N__13071));
    InMux I__1636 (
            .O(N__13079),
            .I(N__13066));
    InMux I__1635 (
            .O(N__13078),
            .I(N__13066));
    InMux I__1634 (
            .O(N__13077),
            .I(N__13063));
    LocalMux I__1633 (
            .O(N__13074),
            .I(N__13060));
    Span4Mux_h I__1632 (
            .O(N__13071),
            .I(N__13057));
    LocalMux I__1631 (
            .O(N__13066),
            .I(\uu2.l_countZ0Z_0 ));
    LocalMux I__1630 (
            .O(N__13063),
            .I(\uu2.l_countZ0Z_0 ));
    Odrv4 I__1629 (
            .O(N__13060),
            .I(\uu2.l_countZ0Z_0 ));
    Odrv4 I__1628 (
            .O(N__13057),
            .I(\uu2.l_countZ0Z_0 ));
    CascadeMux I__1627 (
            .O(N__13048),
            .I(N__13045));
    InMux I__1626 (
            .O(N__13045),
            .I(N__13039));
    InMux I__1625 (
            .O(N__13044),
            .I(N__13039));
    LocalMux I__1624 (
            .O(N__13039),
            .I(N__13036));
    Span4Mux_s3_h I__1623 (
            .O(N__13036),
            .I(N__13033));
    Odrv4 I__1622 (
            .O(N__13033),
            .I(\uu2.un284_ci ));
    CascadeMux I__1621 (
            .O(N__13030),
            .I(\Lab_UT.dictrl.N_9_cascade_ ));
    CascadeMux I__1620 (
            .O(N__13027),
            .I(\Lab_UT.dictrl.N_21_1_cascade_ ));
    InMux I__1619 (
            .O(N__13024),
            .I(N__13018));
    InMux I__1618 (
            .O(N__13023),
            .I(N__13018));
    LocalMux I__1617 (
            .O(N__13018),
            .I(N__13015));
    Odrv4 I__1616 (
            .O(N__13015),
            .I(\uu2.w_data_displaying_2_i_a2_i_a3_1_0 ));
    InMux I__1615 (
            .O(N__13012),
            .I(N__13008));
    InMux I__1614 (
            .O(N__13011),
            .I(N__13004));
    LocalMux I__1613 (
            .O(N__13008),
            .I(N__13001));
    InMux I__1612 (
            .O(N__13007),
            .I(N__12998));
    LocalMux I__1611 (
            .O(N__13004),
            .I(N__12995));
    Span4Mux_v I__1610 (
            .O(N__13001),
            .I(N__12990));
    LocalMux I__1609 (
            .O(N__12998),
            .I(N__12990));
    Span4Mux_h I__1608 (
            .O(N__12995),
            .I(N__12978));
    Span4Mux_v I__1607 (
            .O(N__12990),
            .I(N__12975));
    InMux I__1606 (
            .O(N__12989),
            .I(N__12968));
    InMux I__1605 (
            .O(N__12988),
            .I(N__12968));
    InMux I__1604 (
            .O(N__12987),
            .I(N__12968));
    InMux I__1603 (
            .O(N__12986),
            .I(N__12963));
    InMux I__1602 (
            .O(N__12985),
            .I(N__12963));
    InMux I__1601 (
            .O(N__12984),
            .I(N__12954));
    InMux I__1600 (
            .O(N__12983),
            .I(N__12954));
    InMux I__1599 (
            .O(N__12982),
            .I(N__12954));
    InMux I__1598 (
            .O(N__12981),
            .I(N__12954));
    Span4Mux_v I__1597 (
            .O(N__12978),
            .I(N__12951));
    Odrv4 I__1596 (
            .O(N__12975),
            .I(\uu0.un4_l_count_0 ));
    LocalMux I__1595 (
            .O(N__12968),
            .I(\uu0.un4_l_count_0 ));
    LocalMux I__1594 (
            .O(N__12963),
            .I(\uu0.un4_l_count_0 ));
    LocalMux I__1593 (
            .O(N__12954),
            .I(\uu0.un4_l_count_0 ));
    Odrv4 I__1592 (
            .O(N__12951),
            .I(\uu0.un4_l_count_0 ));
    InMux I__1591 (
            .O(N__12940),
            .I(N__12935));
    InMux I__1590 (
            .O(N__12939),
            .I(N__12932));
    InMux I__1589 (
            .O(N__12938),
            .I(N__12929));
    LocalMux I__1588 (
            .O(N__12935),
            .I(N__12926));
    LocalMux I__1587 (
            .O(N__12932),
            .I(\uu2.un1_l_count_2_0 ));
    LocalMux I__1586 (
            .O(N__12929),
            .I(\uu2.un1_l_count_2_0 ));
    Odrv4 I__1585 (
            .O(N__12926),
            .I(\uu2.un1_l_count_2_0 ));
    InMux I__1584 (
            .O(N__12919),
            .I(N__12916));
    LocalMux I__1583 (
            .O(N__12916),
            .I(N__12912));
    InMux I__1582 (
            .O(N__12915),
            .I(N__12909));
    Span4Mux_h I__1581 (
            .O(N__12912),
            .I(N__12906));
    LocalMux I__1580 (
            .O(N__12909),
            .I(N__12903));
    Span4Mux_v I__1579 (
            .O(N__12906),
            .I(N__12900));
    Span4Mux_h I__1578 (
            .O(N__12903),
            .I(N__12897));
    Odrv4 I__1577 (
            .O(N__12900),
            .I(\uu0.delay_lineZ0Z_0 ));
    Odrv4 I__1576 (
            .O(N__12897),
            .I(\uu0.delay_lineZ0Z_0 ));
    InMux I__1575 (
            .O(N__12892),
            .I(N__12889));
    LocalMux I__1574 (
            .O(N__12889),
            .I(N__12886));
    Odrv12 I__1573 (
            .O(N__12886),
            .I(\uu0.delay_lineZ0Z_1 ));
    InMux I__1572 (
            .O(N__12883),
            .I(N__12880));
    LocalMux I__1571 (
            .O(N__12880),
            .I(\uu2.bitmap_pmux_sn_i7_mux_0 ));
    CascadeMux I__1570 (
            .O(N__12877),
            .I(\uu2.bitmap_pmux_29_0_cascade_ ));
    CascadeMux I__1569 (
            .O(N__12874),
            .I(N__12871));
    InMux I__1568 (
            .O(N__12871),
            .I(N__12865));
    InMux I__1567 (
            .O(N__12870),
            .I(N__12865));
    LocalMux I__1566 (
            .O(N__12865),
            .I(\uu2.bitmap_pmux ));
    InMux I__1565 (
            .O(N__12862),
            .I(N__12859));
    LocalMux I__1564 (
            .O(N__12859),
            .I(\uu2.bitmap_pmux_sn_N_36 ));
    InMux I__1563 (
            .O(N__12856),
            .I(N__12853));
    LocalMux I__1562 (
            .O(N__12853),
            .I(N__12850));
    Span4Mux_h I__1561 (
            .O(N__12850),
            .I(N__12847));
    Odrv4 I__1560 (
            .O(N__12847),
            .I(vbuf_tx_data_6));
    InMux I__1559 (
            .O(N__12844),
            .I(N__12841));
    LocalMux I__1558 (
            .O(N__12841),
            .I(N__12838));
    Span4Mux_v I__1557 (
            .O(N__12838),
            .I(N__12835));
    Odrv4 I__1556 (
            .O(N__12835),
            .I(\buart.Z_tx.shifterZ0Z_7 ));
    CascadeMux I__1555 (
            .O(N__12832),
            .I(N__12827));
    InMux I__1554 (
            .O(N__12831),
            .I(N__12820));
    InMux I__1553 (
            .O(N__12830),
            .I(N__12820));
    InMux I__1552 (
            .O(N__12827),
            .I(N__12808));
    InMux I__1551 (
            .O(N__12826),
            .I(N__12803));
    InMux I__1550 (
            .O(N__12825),
            .I(N__12803));
    LocalMux I__1549 (
            .O(N__12820),
            .I(N__12800));
    InMux I__1548 (
            .O(N__12819),
            .I(N__12781));
    InMux I__1547 (
            .O(N__12818),
            .I(N__12781));
    InMux I__1546 (
            .O(N__12817),
            .I(N__12781));
    InMux I__1545 (
            .O(N__12816),
            .I(N__12781));
    InMux I__1544 (
            .O(N__12815),
            .I(N__12781));
    InMux I__1543 (
            .O(N__12814),
            .I(N__12781));
    InMux I__1542 (
            .O(N__12813),
            .I(N__12781));
    InMux I__1541 (
            .O(N__12812),
            .I(N__12781));
    InMux I__1540 (
            .O(N__12811),
            .I(N__12778));
    LocalMux I__1539 (
            .O(N__12808),
            .I(N__12771));
    LocalMux I__1538 (
            .O(N__12803),
            .I(N__12771));
    Span4Mux_h I__1537 (
            .O(N__12800),
            .I(N__12771));
    InMux I__1536 (
            .O(N__12799),
            .I(N__12766));
    InMux I__1535 (
            .O(N__12798),
            .I(N__12766));
    LocalMux I__1534 (
            .O(N__12781),
            .I(vbuf_tx_data_rdy));
    LocalMux I__1533 (
            .O(N__12778),
            .I(vbuf_tx_data_rdy));
    Odrv4 I__1532 (
            .O(N__12771),
            .I(vbuf_tx_data_rdy));
    LocalMux I__1531 (
            .O(N__12766),
            .I(vbuf_tx_data_rdy));
    InMux I__1530 (
            .O(N__12757),
            .I(N__12754));
    LocalMux I__1529 (
            .O(N__12754),
            .I(N__12751));
    Span4Mux_v I__1528 (
            .O(N__12751),
            .I(N__12748));
    Odrv4 I__1527 (
            .O(N__12748),
            .I(vbuf_tx_data_7));
    CascadeMux I__1526 (
            .O(N__12745),
            .I(N__12742));
    InMux I__1525 (
            .O(N__12742),
            .I(N__12739));
    LocalMux I__1524 (
            .O(N__12739),
            .I(\buart.Z_tx.shifterZ0Z_8 ));
    CEMux I__1523 (
            .O(N__12736),
            .I(N__12733));
    LocalMux I__1522 (
            .O(N__12733),
            .I(N__12730));
    Span4Mux_h I__1521 (
            .O(N__12730),
            .I(N__12726));
    CEMux I__1520 (
            .O(N__12729),
            .I(N__12723));
    Span4Mux_s0_h I__1519 (
            .O(N__12726),
            .I(N__12720));
    LocalMux I__1518 (
            .O(N__12723),
            .I(N__12717));
    Odrv4 I__1517 (
            .O(N__12720),
            .I(\buart.Z_tx.un1_uart_wr_i_0_i ));
    Odrv4 I__1516 (
            .O(N__12717),
            .I(\buart.Z_tx.un1_uart_wr_i_0_i ));
    IoInMux I__1515 (
            .O(N__12712),
            .I(N__12709));
    LocalMux I__1514 (
            .O(N__12709),
            .I(N__12706));
    Span4Mux_s3_h I__1513 (
            .O(N__12706),
            .I(N__12703));
    Odrv4 I__1512 (
            .O(N__12703),
            .I(\uu0.un11_l_count_i ));
    CascadeMux I__1511 (
            .O(N__12700),
            .I(N__12697));
    InMux I__1510 (
            .O(N__12697),
            .I(N__12694));
    LocalMux I__1509 (
            .O(N__12694),
            .I(N__12691));
    Span4Mux_s3_v I__1508 (
            .O(N__12691),
            .I(N__12688));
    Odrv4 I__1507 (
            .O(N__12688),
            .I(\uu2.mem0.w_addr_7 ));
    CascadeMux I__1506 (
            .O(N__12685),
            .I(N__12682));
    InMux I__1505 (
            .O(N__12682),
            .I(N__12679));
    LocalMux I__1504 (
            .O(N__12679),
            .I(N__12676));
    Span4Mux_v I__1503 (
            .O(N__12676),
            .I(N__12673));
    Odrv4 I__1502 (
            .O(N__12673),
            .I(\uu2.mem0.w_addr_1 ));
    CascadeMux I__1501 (
            .O(N__12670),
            .I(\uu2.N_51_cascade_ ));
    InMux I__1500 (
            .O(N__12667),
            .I(N__12661));
    InMux I__1499 (
            .O(N__12666),
            .I(N__12661));
    LocalMux I__1498 (
            .O(N__12661),
            .I(\uu2.N_34 ));
    CascadeMux I__1497 (
            .O(N__12658),
            .I(\uu2.N_34_cascade_ ));
    InMux I__1496 (
            .O(N__12655),
            .I(N__12652));
    LocalMux I__1495 (
            .O(N__12652),
            .I(\uu2.mem0.w_data_0 ));
    CascadeMux I__1494 (
            .O(N__12649),
            .I(\uu2.bitmap_pmux_sn_m15_0_ns_1_cascade_ ));
    InMux I__1493 (
            .O(N__12646),
            .I(N__12643));
    LocalMux I__1492 (
            .O(N__12643),
            .I(\uu2.bitmap_pmux_sn_N_65 ));
    CascadeMux I__1491 (
            .O(N__12640),
            .I(\uu2.bitmap_pmux_sn_m24_0_ns_1_cascade_ ));
    CascadeMux I__1490 (
            .O(N__12637),
            .I(\uu2.bitmap_pmux_sn_i5_mux_cascade_ ));
    CascadeMux I__1489 (
            .O(N__12634),
            .I(N__12631));
    InMux I__1488 (
            .O(N__12631),
            .I(N__12628));
    LocalMux I__1487 (
            .O(N__12628),
            .I(\uu2.mem0.w_addr_8 ));
    InMux I__1486 (
            .O(N__12625),
            .I(N__12622));
    LocalMux I__1485 (
            .O(N__12622),
            .I(N__12619));
    Span4Mux_h I__1484 (
            .O(N__12619),
            .I(N__12616));
    Odrv4 I__1483 (
            .O(N__12616),
            .I(\uu2.vram_rd_clk_detZ0Z_1 ));
    InMux I__1482 (
            .O(N__12613),
            .I(N__12610));
    LocalMux I__1481 (
            .O(N__12610),
            .I(N__12606));
    InMux I__1480 (
            .O(N__12609),
            .I(N__12603));
    Span4Mux_h I__1479 (
            .O(N__12606),
            .I(N__12600));
    LocalMux I__1478 (
            .O(N__12603),
            .I(\uu2.vram_rd_clk_detZ0Z_0 ));
    Odrv4 I__1477 (
            .O(N__12600),
            .I(\uu2.vram_rd_clk_detZ0Z_0 ));
    CEMux I__1476 (
            .O(N__12595),
            .I(N__12592));
    LocalMux I__1475 (
            .O(N__12592),
            .I(N__12589));
    Span4Mux_v I__1474 (
            .O(N__12589),
            .I(N__12586));
    Span4Mux_s1_h I__1473 (
            .O(N__12586),
            .I(N__12583));
    Odrv4 I__1472 (
            .O(N__12583),
            .I(\uu2.vram_rd_clk_det_RNI95711Z0Z_1 ));
    InMux I__1471 (
            .O(N__12580),
            .I(N__12577));
    LocalMux I__1470 (
            .O(N__12577),
            .I(\uu2.mem0.w_data_4 ));
    InMux I__1469 (
            .O(N__12574),
            .I(N__12571));
    LocalMux I__1468 (
            .O(N__12571),
            .I(\uu2.mem0.w_data_5 ));
    InMux I__1467 (
            .O(N__12568),
            .I(N__12565));
    LocalMux I__1466 (
            .O(N__12565),
            .I(\uu2.N_37 ));
    CascadeMux I__1465 (
            .O(N__12562),
            .I(\uu2.N_37_cascade_ ));
    InMux I__1464 (
            .O(N__12559),
            .I(N__12556));
    LocalMux I__1463 (
            .O(N__12556),
            .I(\uu2.mem0.w_data_3 ));
    InMux I__1462 (
            .O(N__12553),
            .I(N__12550));
    LocalMux I__1461 (
            .O(N__12550),
            .I(\uu2.mem0.w_data_1 ));
    InMux I__1460 (
            .O(N__12547),
            .I(N__12544));
    LocalMux I__1459 (
            .O(N__12544),
            .I(\Lab_UT.dictrl.G_19_0_a7_3_2 ));
    InMux I__1458 (
            .O(N__12541),
            .I(N__12538));
    LocalMux I__1457 (
            .O(N__12538),
            .I(G_19_0_a7_4_8));
    InMux I__1456 (
            .O(N__12535),
            .I(N__12532));
    LocalMux I__1455 (
            .O(N__12532),
            .I(G_19_0_a7_4_1));
    CascadeMux I__1454 (
            .O(N__12529),
            .I(N__12526));
    InMux I__1453 (
            .O(N__12526),
            .I(N__12514));
    InMux I__1452 (
            .O(N__12525),
            .I(N__12514));
    InMux I__1451 (
            .O(N__12524),
            .I(N__12514));
    InMux I__1450 (
            .O(N__12523),
            .I(N__12514));
    LocalMux I__1449 (
            .O(N__12514),
            .I(N__12509));
    InMux I__1448 (
            .O(N__12513),
            .I(N__12506));
    InMux I__1447 (
            .O(N__12512),
            .I(N__12503));
    Span4Mux_v I__1446 (
            .O(N__12509),
            .I(N__12498));
    LocalMux I__1445 (
            .O(N__12506),
            .I(N__12498));
    LocalMux I__1444 (
            .O(N__12503),
            .I(\uu0.l_precountZ0Z_0 ));
    Odrv4 I__1443 (
            .O(N__12498),
            .I(\uu0.l_precountZ0Z_0 ));
    InMux I__1442 (
            .O(N__12493),
            .I(N__12490));
    LocalMux I__1441 (
            .O(N__12490),
            .I(N__12487));
    Span4Mux_s1_v I__1440 (
            .O(N__12487),
            .I(N__12484));
    Odrv4 I__1439 (
            .O(N__12484),
            .I(\uu0.un99_ci_0 ));
    InMux I__1438 (
            .O(N__12481),
            .I(N__12475));
    InMux I__1437 (
            .O(N__12480),
            .I(N__12475));
    LocalMux I__1436 (
            .O(N__12475),
            .I(N__12470));
    InMux I__1435 (
            .O(N__12474),
            .I(N__12467));
    InMux I__1434 (
            .O(N__12473),
            .I(N__12464));
    Span4Mux_h I__1433 (
            .O(N__12470),
            .I(N__12461));
    LocalMux I__1432 (
            .O(N__12467),
            .I(N__12458));
    LocalMux I__1431 (
            .O(N__12464),
            .I(\uu0.l_countZ0Z_4 ));
    Odrv4 I__1430 (
            .O(N__12461),
            .I(\uu0.l_countZ0Z_4 ));
    Odrv4 I__1429 (
            .O(N__12458),
            .I(\uu0.l_countZ0Z_4 ));
    InMux I__1428 (
            .O(N__12451),
            .I(N__12446));
    InMux I__1427 (
            .O(N__12450),
            .I(N__12441));
    InMux I__1426 (
            .O(N__12449),
            .I(N__12441));
    LocalMux I__1425 (
            .O(N__12446),
            .I(N__12438));
    LocalMux I__1424 (
            .O(N__12441),
            .I(\uu0.l_countZ0Z_5 ));
    Odrv4 I__1423 (
            .O(N__12438),
            .I(\uu0.l_countZ0Z_5 ));
    CascadeMux I__1422 (
            .O(N__12433),
            .I(N__12430));
    InMux I__1421 (
            .O(N__12430),
            .I(N__12427));
    LocalMux I__1420 (
            .O(N__12427),
            .I(N__12423));
    InMux I__1419 (
            .O(N__12426),
            .I(N__12420));
    Span4Mux_h I__1418 (
            .O(N__12423),
            .I(N__12417));
    LocalMux I__1417 (
            .O(N__12420),
            .I(\uu0.un88_ci_3 ));
    Odrv4 I__1416 (
            .O(N__12417),
            .I(\uu0.un88_ci_3 ));
    InMux I__1415 (
            .O(N__12412),
            .I(N__12406));
    InMux I__1414 (
            .O(N__12411),
            .I(N__12406));
    LocalMux I__1413 (
            .O(N__12406),
            .I(N__12403));
    Span4Mux_v I__1412 (
            .O(N__12403),
            .I(N__12397));
    InMux I__1411 (
            .O(N__12402),
            .I(N__12394));
    InMux I__1410 (
            .O(N__12401),
            .I(N__12389));
    InMux I__1409 (
            .O(N__12400),
            .I(N__12389));
    Odrv4 I__1408 (
            .O(N__12397),
            .I(\uu0.un66_ci ));
    LocalMux I__1407 (
            .O(N__12394),
            .I(\uu0.un66_ci ));
    LocalMux I__1406 (
            .O(N__12389),
            .I(\uu0.un66_ci ));
    CascadeMux I__1405 (
            .O(N__12382),
            .I(\uu0.un88_ci_3_cascade_ ));
    InMux I__1404 (
            .O(N__12379),
            .I(N__12376));
    LocalMux I__1403 (
            .O(N__12376),
            .I(N__12370));
    InMux I__1402 (
            .O(N__12375),
            .I(N__12367));
    InMux I__1401 (
            .O(N__12374),
            .I(N__12364));
    InMux I__1400 (
            .O(N__12373),
            .I(N__12361));
    Span4Mux_s3_h I__1399 (
            .O(N__12370),
            .I(N__12358));
    LocalMux I__1398 (
            .O(N__12367),
            .I(N__12355));
    LocalMux I__1397 (
            .O(N__12364),
            .I(\uu0.l_countZ0Z_6 ));
    LocalMux I__1396 (
            .O(N__12361),
            .I(\uu0.l_countZ0Z_6 ));
    Odrv4 I__1395 (
            .O(N__12358),
            .I(\uu0.l_countZ0Z_6 ));
    Odrv4 I__1394 (
            .O(N__12355),
            .I(\uu0.l_countZ0Z_6 ));
    CEMux I__1393 (
            .O(N__12346),
            .I(N__12331));
    CEMux I__1392 (
            .O(N__12345),
            .I(N__12331));
    CEMux I__1391 (
            .O(N__12344),
            .I(N__12331));
    CEMux I__1390 (
            .O(N__12343),
            .I(N__12331));
    CEMux I__1389 (
            .O(N__12342),
            .I(N__12331));
    GlobalMux I__1388 (
            .O(N__12331),
            .I(N__12328));
    gio2CtrlBuf I__1387 (
            .O(N__12328),
            .I(\uu0.un11_l_count_i_g ));
    InMux I__1386 (
            .O(N__12325),
            .I(N__12322));
    LocalMux I__1385 (
            .O(N__12322),
            .I(\Lab_UT.dictrl.N_5_0_0 ));
    CascadeMux I__1384 (
            .O(N__12319),
            .I(\Lab_UT.dictrl.g0_4_0_cascade_ ));
    CascadeMux I__1383 (
            .O(N__12316),
            .I(\Lab_UT.dictrl.N_8_0_0_cascade_ ));
    InMux I__1382 (
            .O(N__12313),
            .I(N__12310));
    LocalMux I__1381 (
            .O(N__12310),
            .I(\Lab_UT.dictrl.N_4 ));
    InMux I__1380 (
            .O(N__12307),
            .I(N__12304));
    LocalMux I__1379 (
            .O(N__12304),
            .I(\Lab_UT.dictrl.currState_i_5_2 ));
    CascadeMux I__1378 (
            .O(N__12301),
            .I(\Lab_UT.dictrl.G_19_0_a7_4_10_cascade_ ));
    CascadeMux I__1377 (
            .O(N__12298),
            .I(\Lab_UT.dictrl.N_21_cascade_ ));
    InMux I__1376 (
            .O(N__12295),
            .I(N__12292));
    LocalMux I__1375 (
            .O(N__12292),
            .I(N__12289));
    Odrv12 I__1374 (
            .O(N__12289),
            .I(\Lab_UT.dictrl.G_19_0_a7_2_0 ));
    InMux I__1373 (
            .O(N__12286),
            .I(N__12283));
    LocalMux I__1372 (
            .O(N__12283),
            .I(\Lab_UT.dictrl.G_19_0_0 ));
    CascadeMux I__1371 (
            .O(N__12280),
            .I(\Lab_UT.dictrl.i8_mux_0_0_cascade_ ));
    InMux I__1370 (
            .O(N__12277),
            .I(N__12274));
    LocalMux I__1369 (
            .O(N__12274),
            .I(\Lab_UT.dictrl.i7_mux_0 ));
    InMux I__1368 (
            .O(N__12271),
            .I(N__12268));
    LocalMux I__1367 (
            .O(N__12268),
            .I(\Lab_UT.dictrl.N_12 ));
    InMux I__1366 (
            .O(N__12265),
            .I(N__12262));
    LocalMux I__1365 (
            .O(N__12262),
            .I(N__12259));
    Odrv4 I__1364 (
            .O(N__12259),
            .I(\Lab_UT.dictrl.G_30_0_a7_2 ));
    CascadeMux I__1363 (
            .O(N__12256),
            .I(\Lab_UT.dictrl.N_11_0_cascade_ ));
    CascadeMux I__1362 (
            .O(N__12253),
            .I(N__12250));
    InMux I__1361 (
            .O(N__12250),
            .I(N__12247));
    LocalMux I__1360 (
            .O(N__12247),
            .I(\Lab_UT.dictrl.G_30_0_a7_4_1 ));
    InMux I__1359 (
            .O(N__12244),
            .I(N__12241));
    LocalMux I__1358 (
            .O(N__12241),
            .I(\Lab_UT.dictrl.G_30_0_a7_1_2 ));
    CascadeMux I__1357 (
            .O(N__12238),
            .I(\Lab_UT.dictrl.N_31_0_cascade_ ));
    InMux I__1356 (
            .O(N__12235),
            .I(N__12232));
    LocalMux I__1355 (
            .O(N__12232),
            .I(\Lab_UT.dictrl.N_23_1 ));
    CascadeMux I__1354 (
            .O(N__12229),
            .I(\Lab_UT.dictrl.G_30_0_2_cascade_ ));
    CascadeMux I__1353 (
            .O(N__12226),
            .I(\Lab_UT.dictrl.nextStateZ0Z_1_cascade_ ));
    CascadeMux I__1352 (
            .O(N__12223),
            .I(\Lab_UT.dictrl.G_30_0_a7_2_0_cascade_ ));
    InMux I__1351 (
            .O(N__12220),
            .I(N__12217));
    LocalMux I__1350 (
            .O(N__12217),
            .I(\Lab_UT.dictrl.G_30_0_0 ));
    InMux I__1349 (
            .O(N__12214),
            .I(N__12211));
    LocalMux I__1348 (
            .O(N__12211),
            .I(\Lab_UT.dictrl.G_30_0_a7_0_0 ));
    InMux I__1347 (
            .O(N__12208),
            .I(N__12205));
    LocalMux I__1346 (
            .O(N__12205),
            .I(\Lab_UT.dictrl.N_30_0 ));
    InMux I__1345 (
            .O(N__12202),
            .I(N__12187));
    InMux I__1344 (
            .O(N__12201),
            .I(N__12187));
    InMux I__1343 (
            .O(N__12200),
            .I(N__12187));
    InMux I__1342 (
            .O(N__12199),
            .I(N__12187));
    InMux I__1341 (
            .O(N__12198),
            .I(N__12187));
    LocalMux I__1340 (
            .O(N__12187),
            .I(\uu2.l_countZ0Z_6 ));
    CascadeMux I__1339 (
            .O(N__12184),
            .I(N__12178));
    InMux I__1338 (
            .O(N__12183),
            .I(N__12172));
    InMux I__1337 (
            .O(N__12182),
            .I(N__12172));
    InMux I__1336 (
            .O(N__12181),
            .I(N__12165));
    InMux I__1335 (
            .O(N__12178),
            .I(N__12165));
    InMux I__1334 (
            .O(N__12177),
            .I(N__12165));
    LocalMux I__1333 (
            .O(N__12172),
            .I(\uu2.l_countZ0Z_4 ));
    LocalMux I__1332 (
            .O(N__12165),
            .I(\uu2.l_countZ0Z_4 ));
    CascadeMux I__1331 (
            .O(N__12160),
            .I(N__12155));
    InMux I__1330 (
            .O(N__12159),
            .I(N__12148));
    InMux I__1329 (
            .O(N__12158),
            .I(N__12148));
    InMux I__1328 (
            .O(N__12155),
            .I(N__12148));
    LocalMux I__1327 (
            .O(N__12148),
            .I(\uu2.l_countZ0Z_9 ));
    InMux I__1326 (
            .O(N__12145),
            .I(N__12142));
    LocalMux I__1325 (
            .O(N__12142),
            .I(\uu2.un1_l_count_2_2 ));
    CascadeMux I__1324 (
            .O(N__12139),
            .I(\Lab_UT.dictrl.N_8_1_cascade_ ));
    CascadeMux I__1323 (
            .O(N__12136),
            .I(\Lab_UT.dictrl.N_20_0_cascade_ ));
    InMux I__1322 (
            .O(N__12133),
            .I(N__12130));
    LocalMux I__1321 (
            .O(N__12130),
            .I(\Lab_UT.dictrl.N_9_1 ));
    InMux I__1320 (
            .O(N__12127),
            .I(N__12112));
    InMux I__1319 (
            .O(N__12126),
            .I(N__12112));
    InMux I__1318 (
            .O(N__12125),
            .I(N__12112));
    InMux I__1317 (
            .O(N__12124),
            .I(N__12112));
    InMux I__1316 (
            .O(N__12123),
            .I(N__12112));
    LocalMux I__1315 (
            .O(N__12112),
            .I(\uu2.l_countZ0Z_2 ));
    InMux I__1314 (
            .O(N__12109),
            .I(N__12100));
    InMux I__1313 (
            .O(N__12108),
            .I(N__12100));
    InMux I__1312 (
            .O(N__12107),
            .I(N__12100));
    LocalMux I__1311 (
            .O(N__12100),
            .I(\uu2.l_countZ0Z_3 ));
    CascadeMux I__1310 (
            .O(N__12097),
            .I(\uu2.un306_ci_cascade_ ));
    CascadeMux I__1309 (
            .O(N__12094),
            .I(\uu2.un350_ci_cascade_ ));
    InMux I__1308 (
            .O(N__12091),
            .I(N__12088));
    LocalMux I__1307 (
            .O(N__12088),
            .I(\uu2.un1_l_count_1_2_0 ));
    InMux I__1306 (
            .O(N__12085),
            .I(N__12082));
    LocalMux I__1305 (
            .O(N__12082),
            .I(\uu2.un350_ci ));
    CascadeMux I__1304 (
            .O(N__12079),
            .I(N__12074));
    InMux I__1303 (
            .O(N__12078),
            .I(N__12071));
    InMux I__1302 (
            .O(N__12077),
            .I(N__12068));
    InMux I__1301 (
            .O(N__12074),
            .I(N__12065));
    LocalMux I__1300 (
            .O(N__12071),
            .I(\uu2.l_countZ0Z_8 ));
    LocalMux I__1299 (
            .O(N__12068),
            .I(\uu2.l_countZ0Z_8 ));
    LocalMux I__1298 (
            .O(N__12065),
            .I(\uu2.l_countZ0Z_8 ));
    InMux I__1297 (
            .O(N__12058),
            .I(N__12053));
    InMux I__1296 (
            .O(N__12057),
            .I(N__12048));
    InMux I__1295 (
            .O(N__12056),
            .I(N__12048));
    LocalMux I__1294 (
            .O(N__12053),
            .I(\uu2.l_countZ0Z_5 ));
    LocalMux I__1293 (
            .O(N__12048),
            .I(\uu2.l_countZ0Z_5 ));
    CascadeMux I__1292 (
            .O(N__12043),
            .I(N__12039));
    CascadeMux I__1291 (
            .O(N__12042),
            .I(N__12036));
    InMux I__1290 (
            .O(N__12039),
            .I(N__12031));
    InMux I__1289 (
            .O(N__12036),
            .I(N__12031));
    LocalMux I__1288 (
            .O(N__12031),
            .I(\uu2.vbuf_count.un328_ci_3 ));
    CascadeMux I__1287 (
            .O(N__12028),
            .I(\uu2.vbuf_count.un328_ci_3_cascade_ ));
    InMux I__1286 (
            .O(N__12025),
            .I(N__12019));
    InMux I__1285 (
            .O(N__12024),
            .I(N__12012));
    InMux I__1284 (
            .O(N__12023),
            .I(N__12012));
    InMux I__1283 (
            .O(N__12022),
            .I(N__12012));
    LocalMux I__1282 (
            .O(N__12019),
            .I(\uu2.un306_ci ));
    LocalMux I__1281 (
            .O(N__12012),
            .I(\uu2.un306_ci ));
    InMux I__1280 (
            .O(N__12007),
            .I(N__12000));
    InMux I__1279 (
            .O(N__12006),
            .I(N__12000));
    InMux I__1278 (
            .O(N__12005),
            .I(N__11997));
    LocalMux I__1277 (
            .O(N__12000),
            .I(\uu2.l_countZ0Z_7 ));
    LocalMux I__1276 (
            .O(N__11997),
            .I(\uu2.l_countZ0Z_7 ));
    InMux I__1275 (
            .O(N__11992),
            .I(N__11989));
    LocalMux I__1274 (
            .O(N__11989),
            .I(vbuf_tx_data_4));
    InMux I__1273 (
            .O(N__11986),
            .I(N__11983));
    LocalMux I__1272 (
            .O(N__11983),
            .I(\buart.Z_tx.shifterZ0Z_5 ));
    InMux I__1271 (
            .O(N__11980),
            .I(N__11977));
    LocalMux I__1270 (
            .O(N__11977),
            .I(vbuf_tx_data_5));
    InMux I__1269 (
            .O(N__11974),
            .I(N__11971));
    LocalMux I__1268 (
            .O(N__11971),
            .I(\buart.Z_tx.shifterZ0Z_6 ));
    CascadeMux I__1267 (
            .O(N__11968),
            .I(\uu2.un1_l_count_1_3_cascade_ ));
    CascadeMux I__1266 (
            .O(N__11965),
            .I(N__11962));
    InMux I__1265 (
            .O(N__11962),
            .I(N__11959));
    LocalMux I__1264 (
            .O(N__11959),
            .I(\uu2.un1_l_count_1_3 ));
    CascadeMux I__1263 (
            .O(N__11956),
            .I(\uu2.un1_l_count_2_0_cascade_ ));
    InMux I__1262 (
            .O(N__11953),
            .I(N__11950));
    LocalMux I__1261 (
            .O(N__11950),
            .I(\uu2.r_data_wire_6 ));
    InMux I__1260 (
            .O(N__11947),
            .I(N__11944));
    LocalMux I__1259 (
            .O(N__11944),
            .I(\uu2.r_data_wire_7 ));
    InMux I__1258 (
            .O(N__11941),
            .I(N__11938));
    LocalMux I__1257 (
            .O(N__11938),
            .I(vbuf_tx_data_0));
    InMux I__1256 (
            .O(N__11935),
            .I(N__11932));
    LocalMux I__1255 (
            .O(N__11932),
            .I(\buart.Z_tx.shifterZ0Z_1 ));
    InMux I__1254 (
            .O(N__11929),
            .I(N__11926));
    LocalMux I__1253 (
            .O(N__11926),
            .I(\buart.Z_tx.shifterZ0Z_0 ));
    IoInMux I__1252 (
            .O(N__11923),
            .I(N__11920));
    LocalMux I__1251 (
            .O(N__11920),
            .I(N__11917));
    Span4Mux_s1_h I__1250 (
            .O(N__11917),
            .I(N__11914));
    Span4Mux_v I__1249 (
            .O(N__11914),
            .I(N__11911));
    Odrv4 I__1248 (
            .O(N__11911),
            .I(o_serial_data_c));
    InMux I__1247 (
            .O(N__11908),
            .I(N__11905));
    LocalMux I__1246 (
            .O(N__11905),
            .I(vbuf_tx_data_1));
    InMux I__1245 (
            .O(N__11902),
            .I(N__11899));
    LocalMux I__1244 (
            .O(N__11899),
            .I(\buart.Z_tx.shifterZ0Z_2 ));
    InMux I__1243 (
            .O(N__11896),
            .I(N__11893));
    LocalMux I__1242 (
            .O(N__11893),
            .I(vbuf_tx_data_2));
    InMux I__1241 (
            .O(N__11890),
            .I(N__11887));
    LocalMux I__1240 (
            .O(N__11887),
            .I(\buart.Z_tx.shifterZ0Z_3 ));
    InMux I__1239 (
            .O(N__11884),
            .I(N__11881));
    LocalMux I__1238 (
            .O(N__11881),
            .I(vbuf_tx_data_3));
    InMux I__1237 (
            .O(N__11878),
            .I(N__11875));
    LocalMux I__1236 (
            .O(N__11875),
            .I(\buart.Z_tx.shifterZ0Z_4 ));
    InMux I__1235 (
            .O(N__11872),
            .I(N__11857));
    InMux I__1234 (
            .O(N__11871),
            .I(N__11857));
    InMux I__1233 (
            .O(N__11870),
            .I(N__11857));
    InMux I__1232 (
            .O(N__11869),
            .I(N__11857));
    InMux I__1231 (
            .O(N__11868),
            .I(N__11857));
    LocalMux I__1230 (
            .O(N__11857),
            .I(\uu0.l_precountZ0Z_1 ));
    CascadeMux I__1229 (
            .O(N__11854),
            .I(N__11849));
    CascadeMux I__1228 (
            .O(N__11853),
            .I(N__11846));
    InMux I__1227 (
            .O(N__11852),
            .I(N__11839));
    InMux I__1226 (
            .O(N__11849),
            .I(N__11839));
    InMux I__1225 (
            .O(N__11846),
            .I(N__11839));
    LocalMux I__1224 (
            .O(N__11839),
            .I(\uu0.l_precountZ0Z_3 ));
    CascadeMux I__1223 (
            .O(N__11836),
            .I(N__11831));
    InMux I__1222 (
            .O(N__11835),
            .I(N__11823));
    InMux I__1221 (
            .O(N__11834),
            .I(N__11823));
    InMux I__1220 (
            .O(N__11831),
            .I(N__11823));
    InMux I__1219 (
            .O(N__11830),
            .I(N__11820));
    LocalMux I__1218 (
            .O(N__11823),
            .I(\uu0.l_countZ0Z_1 ));
    LocalMux I__1217 (
            .O(N__11820),
            .I(\uu0.l_countZ0Z_1 ));
    InMux I__1216 (
            .O(N__11815),
            .I(N__11811));
    InMux I__1215 (
            .O(N__11814),
            .I(N__11808));
    LocalMux I__1214 (
            .O(N__11811),
            .I(\uu0.l_countZ0Z_18 ));
    LocalMux I__1213 (
            .O(N__11808),
            .I(\uu0.l_countZ0Z_18 ));
    InMux I__1212 (
            .O(N__11803),
            .I(N__11798));
    InMux I__1211 (
            .O(N__11802),
            .I(N__11793));
    InMux I__1210 (
            .O(N__11801),
            .I(N__11793));
    LocalMux I__1209 (
            .O(N__11798),
            .I(N__11790));
    LocalMux I__1208 (
            .O(N__11793),
            .I(\uu0.l_countZ0Z_15 ));
    Odrv4 I__1207 (
            .O(N__11790),
            .I(\uu0.l_countZ0Z_15 ));
    CascadeMux I__1206 (
            .O(N__11785),
            .I(\uu0.un4_l_count_11_cascade_ ));
    InMux I__1205 (
            .O(N__11782),
            .I(N__11779));
    LocalMux I__1204 (
            .O(N__11779),
            .I(N__11776));
    Odrv4 I__1203 (
            .O(N__11776),
            .I(\uu0.un4_l_count_16 ));
    InMux I__1202 (
            .O(N__11773),
            .I(N__11770));
    LocalMux I__1201 (
            .O(N__11770),
            .I(\uu2.r_data_wire_0 ));
    InMux I__1200 (
            .O(N__11767),
            .I(N__11764));
    LocalMux I__1199 (
            .O(N__11764),
            .I(\uu2.r_data_wire_1 ));
    InMux I__1198 (
            .O(N__11761),
            .I(N__11758));
    LocalMux I__1197 (
            .O(N__11758),
            .I(\uu2.r_data_wire_2 ));
    InMux I__1196 (
            .O(N__11755),
            .I(N__11752));
    LocalMux I__1195 (
            .O(N__11752),
            .I(\uu2.r_data_wire_3 ));
    InMux I__1194 (
            .O(N__11749),
            .I(N__11746));
    LocalMux I__1193 (
            .O(N__11746),
            .I(\uu2.r_data_wire_4 ));
    InMux I__1192 (
            .O(N__11743),
            .I(N__11740));
    LocalMux I__1191 (
            .O(N__11740),
            .I(\uu2.r_data_wire_5 ));
    CascadeMux I__1190 (
            .O(N__11737),
            .I(N__11729));
    CascadeMux I__1189 (
            .O(N__11736),
            .I(N__11726));
    CascadeMux I__1188 (
            .O(N__11735),
            .I(N__11720));
    CascadeMux I__1187 (
            .O(N__11734),
            .I(N__11717));
    InMux I__1186 (
            .O(N__11733),
            .I(N__11709));
    InMux I__1185 (
            .O(N__11732),
            .I(N__11709));
    InMux I__1184 (
            .O(N__11729),
            .I(N__11709));
    InMux I__1183 (
            .O(N__11726),
            .I(N__11706));
    InMux I__1182 (
            .O(N__11725),
            .I(N__11699));
    InMux I__1181 (
            .O(N__11724),
            .I(N__11699));
    InMux I__1180 (
            .O(N__11723),
            .I(N__11699));
    InMux I__1179 (
            .O(N__11720),
            .I(N__11692));
    InMux I__1178 (
            .O(N__11717),
            .I(N__11692));
    InMux I__1177 (
            .O(N__11716),
            .I(N__11692));
    LocalMux I__1176 (
            .O(N__11709),
            .I(\uu0.un110_ci ));
    LocalMux I__1175 (
            .O(N__11706),
            .I(\uu0.un110_ci ));
    LocalMux I__1174 (
            .O(N__11699),
            .I(\uu0.un110_ci ));
    LocalMux I__1173 (
            .O(N__11692),
            .I(\uu0.un110_ci ));
    InMux I__1172 (
            .O(N__11683),
            .I(N__11676));
    InMux I__1171 (
            .O(N__11682),
            .I(N__11676));
    InMux I__1170 (
            .O(N__11681),
            .I(N__11673));
    LocalMux I__1169 (
            .O(N__11676),
            .I(N__11670));
    LocalMux I__1168 (
            .O(N__11673),
            .I(\uu0.un198_ci_2 ));
    Odrv4 I__1167 (
            .O(N__11670),
            .I(\uu0.un198_ci_2 ));
    CascadeMux I__1166 (
            .O(N__11665),
            .I(\uu0.un110_ci_cascade_ ));
    InMux I__1165 (
            .O(N__11662),
            .I(N__11654));
    InMux I__1164 (
            .O(N__11661),
            .I(N__11654));
    InMux I__1163 (
            .O(N__11660),
            .I(N__11649));
    InMux I__1162 (
            .O(N__11659),
            .I(N__11649));
    LocalMux I__1161 (
            .O(N__11654),
            .I(\uu0.l_countZ0Z_16 ));
    LocalMux I__1160 (
            .O(N__11649),
            .I(\uu0.l_countZ0Z_16 ));
    CascadeMux I__1159 (
            .O(N__11644),
            .I(\uu0.un220_ci_cascade_ ));
    InMux I__1158 (
            .O(N__11641),
            .I(N__11630));
    InMux I__1157 (
            .O(N__11640),
            .I(N__11630));
    InMux I__1156 (
            .O(N__11639),
            .I(N__11630));
    InMux I__1155 (
            .O(N__11638),
            .I(N__11625));
    InMux I__1154 (
            .O(N__11637),
            .I(N__11625));
    LocalMux I__1153 (
            .O(N__11630),
            .I(\uu0.l_countZ0Z_9 ));
    LocalMux I__1152 (
            .O(N__11625),
            .I(\uu0.l_countZ0Z_9 ));
    CascadeMux I__1151 (
            .O(N__11620),
            .I(N__11617));
    InMux I__1150 (
            .O(N__11617),
            .I(N__11608));
    InMux I__1149 (
            .O(N__11616),
            .I(N__11608));
    InMux I__1148 (
            .O(N__11615),
            .I(N__11608));
    LocalMux I__1147 (
            .O(N__11608),
            .I(\uu0.l_countZ0Z_7 ));
    CascadeMux I__1146 (
            .O(N__11605),
            .I(N__11600));
    InMux I__1145 (
            .O(N__11604),
            .I(N__11593));
    InMux I__1144 (
            .O(N__11603),
            .I(N__11593));
    InMux I__1143 (
            .O(N__11600),
            .I(N__11593));
    LocalMux I__1142 (
            .O(N__11593),
            .I(\uu0.l_countZ0Z_17 ));
    InMux I__1141 (
            .O(N__11590),
            .I(N__11583));
    InMux I__1140 (
            .O(N__11589),
            .I(N__11583));
    InMux I__1139 (
            .O(N__11588),
            .I(N__11580));
    LocalMux I__1138 (
            .O(N__11583),
            .I(\uu0.l_countZ0Z_3 ));
    LocalMux I__1137 (
            .O(N__11580),
            .I(\uu0.l_countZ0Z_3 ));
    InMux I__1136 (
            .O(N__11575),
            .I(N__11572));
    LocalMux I__1135 (
            .O(N__11572),
            .I(\uu0.un4_l_count_12 ));
    InMux I__1134 (
            .O(N__11569),
            .I(N__11566));
    LocalMux I__1133 (
            .O(N__11566),
            .I(N__11560));
    InMux I__1132 (
            .O(N__11565),
            .I(N__11557));
    CascadeMux I__1131 (
            .O(N__11564),
            .I(N__11554));
    CascadeMux I__1130 (
            .O(N__11563),
            .I(N__11551));
    Span4Mux_s2_v I__1129 (
            .O(N__11560),
            .I(N__11547));
    LocalMux I__1128 (
            .O(N__11557),
            .I(N__11544));
    InMux I__1127 (
            .O(N__11554),
            .I(N__11537));
    InMux I__1126 (
            .O(N__11551),
            .I(N__11537));
    InMux I__1125 (
            .O(N__11550),
            .I(N__11537));
    Odrv4 I__1124 (
            .O(N__11547),
            .I(\buart.Z_tx.uart_busy_0_i ));
    Odrv4 I__1123 (
            .O(N__11544),
            .I(\buart.Z_tx.uart_busy_0_i ));
    LocalMux I__1122 (
            .O(N__11537),
            .I(\buart.Z_tx.uart_busy_0_i ));
    InMux I__1121 (
            .O(N__11530),
            .I(N__11527));
    LocalMux I__1120 (
            .O(N__11527),
            .I(N__11520));
    InMux I__1119 (
            .O(N__11526),
            .I(N__11513));
    InMux I__1118 (
            .O(N__11525),
            .I(N__11506));
    InMux I__1117 (
            .O(N__11524),
            .I(N__11506));
    InMux I__1116 (
            .O(N__11523),
            .I(N__11506));
    Span4Mux_s2_v I__1115 (
            .O(N__11520),
            .I(N__11503));
    InMux I__1114 (
            .O(N__11519),
            .I(N__11494));
    InMux I__1113 (
            .O(N__11518),
            .I(N__11494));
    InMux I__1112 (
            .O(N__11517),
            .I(N__11494));
    InMux I__1111 (
            .O(N__11516),
            .I(N__11494));
    LocalMux I__1110 (
            .O(N__11513),
            .I(N__11491));
    LocalMux I__1109 (
            .O(N__11506),
            .I(\buart.Z_tx.ser_clk ));
    Odrv4 I__1108 (
            .O(N__11503),
            .I(\buart.Z_tx.ser_clk ));
    LocalMux I__1107 (
            .O(N__11494),
            .I(\buart.Z_tx.ser_clk ));
    Odrv12 I__1106 (
            .O(N__11491),
            .I(\buart.Z_tx.ser_clk ));
    CascadeMux I__1105 (
            .O(N__11482),
            .I(N__11477));
    InMux I__1104 (
            .O(N__11481),
            .I(N__11474));
    InMux I__1103 (
            .O(N__11480),
            .I(N__11471));
    InMux I__1102 (
            .O(N__11477),
            .I(N__11468));
    LocalMux I__1101 (
            .O(N__11474),
            .I(N__11465));
    LocalMux I__1100 (
            .O(N__11471),
            .I(\buart.Z_tx.bitcountZ0Z_0 ));
    LocalMux I__1099 (
            .O(N__11468),
            .I(\buart.Z_tx.bitcountZ0Z_0 ));
    Odrv4 I__1098 (
            .O(N__11465),
            .I(\buart.Z_tx.bitcountZ0Z_0 ));
    CascadeMux I__1097 (
            .O(N__11458),
            .I(N__11452));
    InMux I__1096 (
            .O(N__11457),
            .I(N__11445));
    InMux I__1095 (
            .O(N__11456),
            .I(N__11445));
    InMux I__1094 (
            .O(N__11455),
            .I(N__11445));
    InMux I__1093 (
            .O(N__11452),
            .I(N__11442));
    LocalMux I__1092 (
            .O(N__11445),
            .I(\uu0.l_precountZ0Z_2 ));
    LocalMux I__1091 (
            .O(N__11442),
            .I(\uu0.l_precountZ0Z_2 ));
    InMux I__1090 (
            .O(N__11437),
            .I(N__11434));
    LocalMux I__1089 (
            .O(N__11434),
            .I(\uu0.un4_l_count_13 ));
    CascadeMux I__1088 (
            .O(N__11431),
            .I(\uu0.un4_l_count_18_cascade_ ));
    CascadeMux I__1087 (
            .O(N__11428),
            .I(\uu0.un4_l_count_0_cascade_ ));
    InMux I__1086 (
            .O(N__11425),
            .I(N__11422));
    LocalMux I__1085 (
            .O(N__11422),
            .I(\uu0.un143_ci_0 ));
    CascadeMux I__1084 (
            .O(N__11419),
            .I(N__11415));
    InMux I__1083 (
            .O(N__11418),
            .I(N__11409));
    InMux I__1082 (
            .O(N__11415),
            .I(N__11409));
    InMux I__1081 (
            .O(N__11414),
            .I(N__11406));
    LocalMux I__1080 (
            .O(N__11409),
            .I(\uu0.l_countZ0Z_11 ));
    LocalMux I__1079 (
            .O(N__11406),
            .I(\uu0.l_countZ0Z_11 ));
    CascadeMux I__1078 (
            .O(N__11401),
            .I(N__11398));
    InMux I__1077 (
            .O(N__11398),
            .I(N__11386));
    InMux I__1076 (
            .O(N__11397),
            .I(N__11386));
    InMux I__1075 (
            .O(N__11396),
            .I(N__11386));
    InMux I__1074 (
            .O(N__11395),
            .I(N__11386));
    LocalMux I__1073 (
            .O(N__11386),
            .I(\uu0.l_countZ0Z_10 ));
    InMux I__1072 (
            .O(N__11383),
            .I(N__11375));
    InMux I__1071 (
            .O(N__11382),
            .I(N__11375));
    InMux I__1070 (
            .O(N__11381),
            .I(N__11370));
    InMux I__1069 (
            .O(N__11380),
            .I(N__11370));
    LocalMux I__1068 (
            .O(N__11375),
            .I(\uu0.un154_ci_9 ));
    LocalMux I__1067 (
            .O(N__11370),
            .I(\uu0.un154_ci_9 ));
    CascadeMux I__1066 (
            .O(N__11365),
            .I(\uu0.un154_ci_9_cascade_ ));
    InMux I__1065 (
            .O(N__11362),
            .I(N__11357));
    InMux I__1064 (
            .O(N__11361),
            .I(N__11352));
    InMux I__1063 (
            .O(N__11360),
            .I(N__11352));
    LocalMux I__1062 (
            .O(N__11357),
            .I(\uu0.un4_l_count_0_8 ));
    LocalMux I__1061 (
            .O(N__11352),
            .I(\uu0.un4_l_count_0_8 ));
    CascadeMux I__1060 (
            .O(N__11347),
            .I(N__11341));
    InMux I__1059 (
            .O(N__11346),
            .I(N__11336));
    InMux I__1058 (
            .O(N__11345),
            .I(N__11336));
    InMux I__1057 (
            .O(N__11344),
            .I(N__11331));
    InMux I__1056 (
            .O(N__11341),
            .I(N__11331));
    LocalMux I__1055 (
            .O(N__11336),
            .I(\uu0.l_countZ0Z_14 ));
    LocalMux I__1054 (
            .O(N__11331),
            .I(\uu0.l_countZ0Z_14 ));
    InMux I__1053 (
            .O(N__11326),
            .I(N__11318));
    InMux I__1052 (
            .O(N__11325),
            .I(N__11313));
    InMux I__1051 (
            .O(N__11324),
            .I(N__11313));
    InMux I__1050 (
            .O(N__11323),
            .I(N__11306));
    InMux I__1049 (
            .O(N__11322),
            .I(N__11306));
    InMux I__1048 (
            .O(N__11321),
            .I(N__11306));
    LocalMux I__1047 (
            .O(N__11318),
            .I(\uu0.l_countZ0Z_8 ));
    LocalMux I__1046 (
            .O(N__11313),
            .I(\uu0.l_countZ0Z_8 ));
    LocalMux I__1045 (
            .O(N__11306),
            .I(\uu0.l_countZ0Z_8 ));
    CascadeMux I__1044 (
            .O(N__11299),
            .I(\Lab_UT.dictrl.currState_0_ret_28_RNOZ0Z_4_cascade_ ));
    InMux I__1043 (
            .O(N__11296),
            .I(N__11293));
    LocalMux I__1042 (
            .O(N__11293),
            .I(\Lab_UT.dictrl.N_1605_0 ));
    InMux I__1041 (
            .O(N__11290),
            .I(N__11287));
    LocalMux I__1040 (
            .O(N__11287),
            .I(\Lab_UT.dictrl.N_5_0 ));
    CascadeMux I__1039 (
            .O(N__11284),
            .I(\Lab_UT.dictrl.g1_0_cascade_ ));
    CascadeMux I__1038 (
            .O(N__11281),
            .I(\Lab_UT.dictrl.g0_i_o4_4_1_cascade_ ));
    CascadeMux I__1037 (
            .O(N__11278),
            .I(\Lab_UT.dictrl.g0_i_o4_4_cascade_ ));
    InMux I__1036 (
            .O(N__11275),
            .I(N__11272));
    LocalMux I__1035 (
            .O(N__11272),
            .I(uart_RXD));
    InMux I__1034 (
            .O(N__11269),
            .I(N__11259));
    InMux I__1033 (
            .O(N__11268),
            .I(N__11259));
    InMux I__1032 (
            .O(N__11267),
            .I(N__11259));
    InMux I__1031 (
            .O(N__11266),
            .I(N__11256));
    LocalMux I__1030 (
            .O(N__11259),
            .I(\uu0.l_countZ0Z_2 ));
    LocalMux I__1029 (
            .O(N__11256),
            .I(\uu0.l_countZ0Z_2 ));
    CascadeMux I__1028 (
            .O(N__11251),
            .I(\uu0.un4_l_count_14_cascade_ ));
    CascadeMux I__1027 (
            .O(N__11248),
            .I(\Lab_UT.dictrl.N_17_1_cascade_ ));
    CascadeMux I__1026 (
            .O(N__11245),
            .I(\Lab_UT.dictrl.g0_i_4_0_cascade_ ));
    InMux I__1025 (
            .O(N__11242),
            .I(N__11239));
    LocalMux I__1024 (
            .O(N__11239),
            .I(\Lab_UT.dictrl.N_19 ));
    CascadeMux I__1023 (
            .O(N__11236),
            .I(N__11233));
    InMux I__1022 (
            .O(N__11233),
            .I(N__11230));
    LocalMux I__1021 (
            .O(N__11230),
            .I(\Lab_UT.dictrl.N_8_2 ));
    CascadeMux I__1020 (
            .O(N__11227),
            .I(\Lab_UT.dictrl.N_8_2_cascade_ ));
    InMux I__1019 (
            .O(N__11224),
            .I(N__11221));
    LocalMux I__1018 (
            .O(N__11221),
            .I(\Lab_UT.dictrl.g0_i_a8_0_1 ));
    InMux I__1017 (
            .O(N__11218),
            .I(N__11215));
    LocalMux I__1016 (
            .O(N__11215),
            .I(\Lab_UT.dictrl.N_1605_1 ));
    InMux I__1015 (
            .O(N__11212),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_2 ));
    InMux I__1014 (
            .O(N__11209),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_3 ));
    InMux I__1013 (
            .O(N__11206),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_4 ));
    InMux I__1012 (
            .O(N__11203),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_5 ));
    CascadeMux I__1011 (
            .O(N__11200),
            .I(N__11197));
    InMux I__1010 (
            .O(N__11197),
            .I(N__11191));
    InMux I__1009 (
            .O(N__11196),
            .I(N__11191));
    LocalMux I__1008 (
            .O(N__11191),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_5 ));
    CascadeMux I__1007 (
            .O(N__11188),
            .I(N__11185));
    InMux I__1006 (
            .O(N__11185),
            .I(N__11179));
    InMux I__1005 (
            .O(N__11184),
            .I(N__11179));
    LocalMux I__1004 (
            .O(N__11179),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_4 ));
    CascadeMux I__1003 (
            .O(N__11176),
            .I(N__11172));
    InMux I__1002 (
            .O(N__11175),
            .I(N__11169));
    InMux I__1001 (
            .O(N__11172),
            .I(N__11166));
    LocalMux I__1000 (
            .O(N__11169),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_6 ));
    LocalMux I__999 (
            .O(N__11166),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_6 ));
    InMux I__998 (
            .O(N__11161),
            .I(N__11155));
    InMux I__997 (
            .O(N__11160),
            .I(N__11155));
    LocalMux I__996 (
            .O(N__11155),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_3 ));
    InMux I__995 (
            .O(N__11152),
            .I(N__11146));
    InMux I__994 (
            .O(N__11151),
            .I(N__11146));
    LocalMux I__993 (
            .O(N__11146),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_2 ));
    CascadeMux I__992 (
            .O(N__11143),
            .I(\buart.Z_tx.Z_baudgen.ser_clk_4_cascade_ ));
    CascadeMux I__991 (
            .O(N__11140),
            .I(N__11136));
    InMux I__990 (
            .O(N__11139),
            .I(N__11132));
    InMux I__989 (
            .O(N__11136),
            .I(N__11127));
    InMux I__988 (
            .O(N__11135),
            .I(N__11127));
    LocalMux I__987 (
            .O(N__11132),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_1 ));
    LocalMux I__986 (
            .O(N__11127),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_1 ));
    InMux I__985 (
            .O(N__11122),
            .I(N__11114));
    InMux I__984 (
            .O(N__11121),
            .I(N__11114));
    InMux I__983 (
            .O(N__11120),
            .I(N__11109));
    InMux I__982 (
            .O(N__11119),
            .I(N__11109));
    LocalMux I__981 (
            .O(N__11114),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_0 ));
    LocalMux I__980 (
            .O(N__11109),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_0 ));
    InMux I__979 (
            .O(N__11104),
            .I(\buart.Z_tx.un1_bitcount_cry_1 ));
    InMux I__978 (
            .O(N__11101),
            .I(\buart.Z_tx.un1_bitcount_cry_2 ));
    InMux I__977 (
            .O(N__11098),
            .I(N__11095));
    LocalMux I__976 (
            .O(N__11095),
            .I(\buart.Z_tx.bitcount_RNIVE1P1Z0Z_3 ));
    InMux I__975 (
            .O(N__11092),
            .I(N__11089));
    LocalMux I__974 (
            .O(N__11089),
            .I(\buart.Z_tx.un1_bitcount_axb_3 ));
    InMux I__973 (
            .O(N__11086),
            .I(N__11083));
    LocalMux I__972 (
            .O(N__11083),
            .I(\buart.Z_tx.un1_bitcount_cry_0_0_c_RNOZ0 ));
    CascadeMux I__971 (
            .O(N__11080),
            .I(N__11077));
    InMux I__970 (
            .O(N__11077),
            .I(N__11073));
    InMux I__969 (
            .O(N__11076),
            .I(N__11070));
    LocalMux I__968 (
            .O(N__11073),
            .I(\buart.Z_tx.bitcountZ0Z_1 ));
    LocalMux I__967 (
            .O(N__11070),
            .I(\buart.Z_tx.bitcountZ0Z_1 ));
    CascadeMux I__966 (
            .O(N__11065),
            .I(N__11061));
    InMux I__965 (
            .O(N__11064),
            .I(N__11058));
    InMux I__964 (
            .O(N__11061),
            .I(N__11055));
    LocalMux I__963 (
            .O(N__11058),
            .I(\buart.Z_tx.bitcountZ0Z_3 ));
    LocalMux I__962 (
            .O(N__11055),
            .I(\buart.Z_tx.bitcountZ0Z_3 ));
    CascadeMux I__961 (
            .O(N__11050),
            .I(N__11047));
    InMux I__960 (
            .O(N__11047),
            .I(N__11043));
    InMux I__959 (
            .O(N__11046),
            .I(N__11040));
    LocalMux I__958 (
            .O(N__11043),
            .I(\buart.Z_tx.bitcountZ0Z_2 ));
    LocalMux I__957 (
            .O(N__11040),
            .I(\buart.Z_tx.bitcountZ0Z_2 ));
    CascadeMux I__956 (
            .O(N__11035),
            .I(\buart.Z_tx.uart_busy_0_i_cascade_ ));
    InMux I__955 (
            .O(N__11032),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_1 ));
    CascadeMux I__954 (
            .O(N__11029),
            .I(N__11024));
    InMux I__953 (
            .O(N__11028),
            .I(N__11011));
    InMux I__952 (
            .O(N__11027),
            .I(N__11011));
    InMux I__951 (
            .O(N__11024),
            .I(N__11011));
    InMux I__950 (
            .O(N__11023),
            .I(N__11011));
    InMux I__949 (
            .O(N__11022),
            .I(N__11011));
    LocalMux I__948 (
            .O(N__11011),
            .I(\uu0.l_countZ0Z_0 ));
    CascadeMux I__947 (
            .O(N__11008),
            .I(N__11005));
    InMux I__946 (
            .O(N__11005),
            .I(N__11002));
    LocalMux I__945 (
            .O(N__11002),
            .I(\uu0.un44_ci ));
    CascadeMux I__944 (
            .O(N__10999),
            .I(\uu0.un44_ci_cascade_ ));
    InMux I__943 (
            .O(N__10996),
            .I(\buart.Z_tx.un1_bitcount_cry_0 ));
    InMux I__942 (
            .O(N__10993),
            .I(N__10990));
    LocalMux I__941 (
            .O(N__10990),
            .I(\buart.Z_tx.bitcount_RNIVE1P1_0Z0Z_3 ));
    CascadeMux I__940 (
            .O(N__10987),
            .I(\uu0.un187_ci_1_cascade_ ));
    InMux I__939 (
            .O(N__10984),
            .I(N__10981));
    LocalMux I__938 (
            .O(N__10981),
            .I(\uu0.un165_ci_0 ));
    CascadeMux I__937 (
            .O(N__10978),
            .I(N__10975));
    InMux I__936 (
            .O(N__10975),
            .I(N__10969));
    InMux I__935 (
            .O(N__10974),
            .I(N__10969));
    LocalMux I__934 (
            .O(N__10969),
            .I(\uu0.l_countZ0Z_13 ));
    InMux I__933 (
            .O(N__10966),
            .I(N__10957));
    InMux I__932 (
            .O(N__10965),
            .I(N__10957));
    InMux I__931 (
            .O(N__10964),
            .I(N__10957));
    LocalMux I__930 (
            .O(N__10957),
            .I(\uu0.l_countZ0Z_12 ));
    CascadeMux I__929 (
            .O(N__10954),
            .I(\uu0.un4_l_count_0_8_cascade_ ));
    IoInMux I__928 (
            .O(N__10951),
            .I(N__10948));
    LocalMux I__927 (
            .O(N__10948),
            .I(N__10945));
    Span12Mux_s9_v I__926 (
            .O(N__10945),
            .I(N__10942));
    Odrv12 I__925 (
            .O(N__10942),
            .I(\latticehx1k_pll_inst.clk ));
    IoInMux I__924 (
            .O(N__10939),
            .I(N__10936));
    LocalMux I__923 (
            .O(N__10936),
            .I(N__10933));
    IoSpan4Mux I__922 (
            .O(N__10933),
            .I(N__10930));
    Odrv4 I__921 (
            .O(N__10930),
            .I(clk_in_c));
    INV \INVuu2.w_addr_user_5C  (
            .O(\INVuu2.w_addr_user_5C_net ),
            .I(N__29465));
    INV \INVuu2.bitmap_93C  (
            .O(\INVuu2.bitmap_93C_net ),
            .I(N__29435));
    INV \INVuu2.w_addr_user_0C  (
            .O(\INVuu2.w_addr_user_0C_net ),
            .I(N__29449));
    INV \INVuu2.bitmap_212C  (
            .O(\INVuu2.bitmap_212C_net ),
            .I(N__29416));
    INV \INVuu2.bitmap_90C  (
            .O(\INVuu2.bitmap_90C_net ),
            .I(N__29425));
    INV \INVuu2.bitmap_308C  (
            .O(\INVuu2.bitmap_308C_net ),
            .I(N__29434));
    INV \INVuu2.w_addr_displaying_8C  (
            .O(\INVuu2.w_addr_displaying_8C_net ),
            .I(N__29440));
    INV \INVuu2.w_addr_user_nesr_3C  (
            .O(\INVuu2.w_addr_user_nesr_3C_net ),
            .I(N__29448));
    INV \INVuu2.bitmap_194C  (
            .O(\INVuu2.bitmap_194C_net ),
            .I(N__29398));
    INV \INVuu2.bitmap_203C  (
            .O(\INVuu2.bitmap_203C_net ),
            .I(N__29404));
    INV \INVuu2.bitmap_87C  (
            .O(\INVuu2.bitmap_87C_net ),
            .I(N__29411));
    INV \INVuu2.w_addr_displaying_nesr_3C  (
            .O(\INVuu2.w_addr_displaying_nesr_3C_net ),
            .I(N__29418));
    INV \INVuu2.bitmap_111C  (
            .O(\INVuu2.bitmap_111C_net ),
            .I(N__29428));
    INV \INVuu2.bitmap_72C  (
            .O(\INVuu2.bitmap_72C_net ),
            .I(N__29415));
    INV \INVuu2.bitmap_197C  (
            .O(\INVuu2.bitmap_197C_net ),
            .I(N__29424));
    INV \INVuu2.bitmap_290C  (
            .O(\INVuu2.bitmap_290C_net ),
            .I(N__29433));
    INV \INVuu2.vram_rd_clk_det_0C  (
            .O(\INVuu2.vram_rd_clk_det_0C_net ),
            .I(N__29446));
    INV \INVuu2.r_data_reg_0C  (
            .O(\INVuu2.r_data_reg_0C_net ),
            .I(N__29460));
    defparam IN_MUX_bfv_1_4_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_4_0_));
    defparam IN_MUX_bfv_1_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_6_0_));
    defparam IN_MUX_bfv_6_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_16_0_));
    defparam IN_MUX_bfv_4_16_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_16_0_));
    defparam IN_MUX_bfv_12_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_9_0_));
    ICE_GB \latticehx1k_pll_inst.latticehx1k_pll_inst_RNIQV8B  (
            .USERSIGNALTOGLOBALBUFFER(N__10951),
            .GLOBALBUFFEROUTPUT(clk_g));
    ICE_GB \buart.Z_rx.bitcount_es_RNIV4M42_0_0  (
            .USERSIGNALTOGLOBALBUFFER(N__15649),
            .GLOBALBUFFEROUTPUT(\buart.Z_rx.sample_g ));
    ICE_GB \Lab_UT.uu0.delay_line_RNII8EF5_0_1  (
            .USERSIGNALTOGLOBALBUFFER(N__19111),
            .GLOBALBUFFEROUTPUT(\Lab_UT.uu0.un11_l_count_i_g ));
    ICE_GB \uu0.delay_line_RNILLLG7_0_1  (
            .USERSIGNALTOGLOBALBUFFER(N__12712),
            .GLOBALBUFFEROUTPUT(\uu0.un11_l_count_i_g ));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    ICE_GB \resetGen.rst_RNI4PQ1  (
            .USERSIGNALTOGLOBALBUFFER(N__24702),
            .GLOBALBUFFEROUTPUT(rst_g));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \uu0.l_count_13_LC_1_1_0 .C_ON=1'b0;
    defparam \uu0.l_count_13_LC_1_1_0 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_13_LC_1_1_0 .LUT_INIT=16'b0001010001010000;
    LogicCell40 \uu0.l_count_13_LC_1_1_0  (
            .in0(N__12982),
            .in1(N__10984),
            .in2(N__10978),
            .in3(N__11732),
            .lcout(\uu0.l_countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29480),
            .ce(N__12343),
            .sr(N__26085));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_1_1_1 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_1_1_1 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_1_1_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_1_1_1  (
            .in0(N__11346),
            .in1(N__11381),
            .in2(_gnd_net_),
            .in3(N__11362),
            .lcout(),
            .ltout(\uu0.un187_ci_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_15_LC_1_1_2 .C_ON=1'b0;
    defparam \uu0.l_count_15_LC_1_1_2 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_15_LC_1_1_2 .LUT_INIT=16'b0001010101000000;
    LogicCell40 \uu0.l_count_15_LC_1_1_2  (
            .in0(N__12983),
            .in1(N__11733),
            .in2(N__10987),
            .in3(N__11802),
            .lcout(\uu0.l_countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29480),
            .ce(N__12343),
            .sr(N__26085));
    defparam \uu0.l_count_12_LC_1_1_3 .C_ON=1'b0;
    defparam \uu0.l_count_12_LC_1_1_3 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_12_LC_1_1_3 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \uu0.l_count_12_LC_1_1_3  (
            .in0(N__11383),
            .in1(N__10966),
            .in2(N__11737),
            .in3(N__12981),
            .lcout(\uu0.l_countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29480),
            .ce(N__12343),
            .sr(N__26085));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_1_1_4 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_1_1_4 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_1_1_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_1_1_4  (
            .in0(N__10965),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11382),
            .lcout(\uu0.un165_ci_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_RNIFAQ9_13_LC_1_1_5 .C_ON=1'b0;
    defparam \uu0.l_count_RNIFAQ9_13_LC_1_1_5 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNIFAQ9_13_LC_1_1_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu0.l_count_RNIFAQ9_13_LC_1_1_5  (
            .in0(_gnd_net_),
            .in1(N__10974),
            .in2(_gnd_net_),
            .in3(N__10964),
            .lcout(\uu0.un4_l_count_0_8 ),
            .ltout(\uu0.un4_l_count_0_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_1_1_6 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_1_1_6 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_1_1_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_1_1_6  (
            .in0(N__11380),
            .in1(N__11801),
            .in2(N__10954),
            .in3(N__11345),
            .lcout(\uu0.un198_ci_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_4_LC_1_1_7 .C_ON=1'b0;
    defparam \uu0.l_count_4_LC_1_1_7 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_4_LC_1_1_7 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \uu0.l_count_4_LC_1_1_7  (
            .in0(N__12402),
            .in1(N__12473),
            .in2(_gnd_net_),
            .in3(N__12984),
            .lcout(\uu0.l_countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29480),
            .ce(N__12343),
            .sr(N__26085));
    defparam \uu0.l_count_RNI2CNU_11_LC_1_2_0 .C_ON=1'b0;
    defparam \uu0.l_count_RNI2CNU_11_LC_1_2_0 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNI2CNU_11_LC_1_2_0 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \uu0.l_count_RNI2CNU_11_LC_1_2_0  (
            .in0(N__11414),
            .in1(N__11659),
            .in2(N__11458),
            .in3(N__11022),
            .lcout(\uu0.un4_l_count_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_3_LC_1_2_1 .C_ON=1'b0;
    defparam \uu0.l_count_3_LC_1_2_1 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_3_LC_1_2_1 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \uu0.l_count_3_LC_1_2_1  (
            .in0(N__11269),
            .in1(N__11590),
            .in2(N__11008),
            .in3(N__12989),
            .lcout(\uu0.l_countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29478),
            .ce(N__12342),
            .sr(N__26083));
    defparam \uu0.l_count_1_LC_1_2_2 .C_ON=1'b0;
    defparam \uu0.l_count_1_LC_1_2_2 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_1_LC_1_2_2 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \uu0.l_count_1_LC_1_2_2  (
            .in0(N__11835),
            .in1(N__11028),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uu0.l_countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29478),
            .ce(N__12342),
            .sr(N__26083));
    defparam \uu0.l_count_0_LC_1_2_3 .C_ON=1'b0;
    defparam \uu0.l_count_0_LC_1_2_3 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_0_LC_1_2_3 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \uu0.l_count_0_LC_1_2_3  (
            .in0(N__11027),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12987),
            .lcout(\uu0.l_countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29478),
            .ce(N__12342),
            .sr(N__26083));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_1_2_4 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_1_2_4 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_1_2_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_1_2_4  (
            .in0(N__11589),
            .in1(N__11267),
            .in2(N__11836),
            .in3(N__11023),
            .lcout(\uu0.un66_ci ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_1_LC_1_2_5 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_1_LC_1_2_5 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_1_LC_1_2_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_1_LC_1_2_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11029),
            .in3(N__11834),
            .lcout(\uu0.un44_ci ),
            .ltout(\uu0.un44_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_2_LC_1_2_6 .C_ON=1'b0;
    defparam \uu0.l_count_2_LC_1_2_6 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_2_LC_1_2_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \uu0.l_count_2_LC_1_2_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10999),
            .in3(N__11268),
            .lcout(\uu0.l_countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29478),
            .ce(N__12342),
            .sr(N__26083));
    defparam \uu0.l_count_16_LC_1_2_7 .C_ON=1'b0;
    defparam \uu0.l_count_16_LC_1_2_7 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_16_LC_1_2_7 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \uu0.l_count_16_LC_1_2_7  (
            .in0(N__11660),
            .in1(N__11681),
            .in2(N__11736),
            .in3(N__12988),
            .lcout(\uu0.l_countZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29478),
            .ce(N__12342),
            .sr(N__26083));
    defparam \buart.Z_tx.bitcount_RNIVE1P1_0_3_LC_1_3_3 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNIVE1P1_0_3_LC_1_3_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNIVE1P1_0_3_LC_1_3_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \buart.Z_tx.bitcount_RNIVE1P1_0_3_LC_1_3_3  (
            .in0(_gnd_net_),
            .in1(N__11565),
            .in2(_gnd_net_),
            .in3(N__11526),
            .lcout(\buart.Z_tx.bitcount_RNIVE1P1_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.un1_bitcount_cry_0_0_c_LC_1_4_0 .C_ON=1'b1;
    defparam \buart.Z_tx.un1_bitcount_cry_0_0_c_LC_1_4_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.un1_bitcount_cry_0_0_c_LC_1_4_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \buart.Z_tx.un1_bitcount_cry_0_0_c_LC_1_4_0  (
            .in0(_gnd_net_),
            .in1(N__11086),
            .in2(N__11482),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_4_0_),
            .carryout(\buart.Z_tx.un1_bitcount_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_1_LC_1_4_1 .C_ON=1'b1;
    defparam \buart.Z_tx.bitcount_1_LC_1_4_1 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.bitcount_1_LC_1_4_1 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \buart.Z_tx.bitcount_1_LC_1_4_1  (
            .in0(N__12825),
            .in1(N__11098),
            .in2(N__11080),
            .in3(N__10996),
            .lcout(\buart.Z_tx.bitcountZ0Z_1 ),
            .ltout(),
            .carryin(\buart.Z_tx.un1_bitcount_cry_0 ),
            .carryout(\buart.Z_tx.un1_bitcount_cry_1 ),
            .clk(N__29468),
            .ce(),
            .sr(N__26079));
    defparam \buart.Z_tx.bitcount_2_LC_1_4_2 .C_ON=1'b1;
    defparam \buart.Z_tx.bitcount_2_LC_1_4_2 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.bitcount_2_LC_1_4_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \buart.Z_tx.bitcount_2_LC_1_4_2  (
            .in0(N__12811),
            .in1(N__10993),
            .in2(N__11050),
            .in3(N__11104),
            .lcout(\buart.Z_tx.bitcountZ0Z_2 ),
            .ltout(),
            .carryin(\buart.Z_tx.un1_bitcount_cry_1 ),
            .carryout(\buart.Z_tx.un1_bitcount_cry_2 ),
            .clk(N__29468),
            .ce(),
            .sr(N__26079));
    defparam \buart.Z_tx.bitcount_3_LC_1_4_3 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_3_LC_1_4_3 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.bitcount_3_LC_1_4_3 .LUT_INIT=16'b1011101111101110;
    LogicCell40 \buart.Z_tx.bitcount_3_LC_1_4_3  (
            .in0(N__12826),
            .in1(N__11092),
            .in2(_gnd_net_),
            .in3(N__11101),
            .lcout(\buart.Z_tx.bitcountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29468),
            .ce(),
            .sr(N__26079));
    defparam \buart.Z_tx.bitcount_RNIVE1P1_3_LC_1_5_0 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNIVE1P1_3_LC_1_5_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNIVE1P1_3_LC_1_5_0 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \buart.Z_tx.bitcount_RNIVE1P1_3_LC_1_5_0  (
            .in0(N__11518),
            .in1(_gnd_net_),
            .in2(N__11563),
            .in3(_gnd_net_),
            .lcout(\buart.Z_tx.bitcount_RNIVE1P1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_data_rdy_LC_1_5_3 .C_ON=1'b0;
    defparam \uu2.r_data_rdy_LC_1_5_3 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_rdy_LC_1_5_3 .LUT_INIT=16'b1111100000001000;
    LogicCell40 \uu2.r_data_rdy_LC_1_5_3  (
            .in0(N__13468),
            .in1(N__13425),
            .in2(N__26158),
            .in3(N__12799),
            .lcout(vbuf_tx_data_rdy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29459),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNO_0_3_LC_1_5_4 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNO_0_3_LC_1_5_4 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNO_0_3_LC_1_5_4 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \buart.Z_tx.bitcount_RNO_0_3_LC_1_5_4  (
            .in0(N__11519),
            .in1(_gnd_net_),
            .in2(N__11564),
            .in3(N__11064),
            .lcout(\buart.Z_tx.un1_bitcount_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.un1_bitcount_cry_0_0_c_RNO_LC_1_5_5 .C_ON=1'b0;
    defparam \buart.Z_tx.un1_bitcount_cry_0_0_c_RNO_LC_1_5_5 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.un1_bitcount_cry_0_0_c_RNO_LC_1_5_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \buart.Z_tx.un1_bitcount_cry_0_0_c_RNO_LC_1_5_5  (
            .in0(_gnd_net_),
            .in1(N__11550),
            .in2(_gnd_net_),
            .in3(N__11517),
            .lcout(\buart.Z_tx.un1_bitcount_cry_0_0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNIQOQA1_3_LC_1_5_6 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNIQOQA1_3_LC_1_5_6 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNIQOQA1_3_LC_1_5_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \buart.Z_tx.bitcount_RNIQOQA1_3_LC_1_5_6  (
            .in0(N__11481),
            .in1(N__11076),
            .in2(N__11065),
            .in3(N__11046),
            .lcout(\buart.Z_tx.uart_busy_0_i ),
            .ltout(\buart.Z_tx.uart_busy_0_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNI22V22_3_LC_1_5_7 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNI22V22_3_LC_1_5_7 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNI22V22_3_LC_1_5_7 .LUT_INIT=16'b1111110011001100;
    LogicCell40 \buart.Z_tx.bitcount_RNI22V22_3_LC_1_5_7  (
            .in0(_gnd_net_),
            .in1(N__12798),
            .in2(N__11035),
            .in3(N__11516),
            .lcout(\buart.Z_tx.un1_uart_wr_i_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_1_6_0 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_1_6_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_1_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_1_6_0  (
            .in0(_gnd_net_),
            .in1(N__11120),
            .in2(N__11140),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_6_0_),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_2_LC_1_6_1 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_2_LC_1_6_1 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_2_LC_1_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_2_LC_1_6_1  (
            .in0(_gnd_net_),
            .in1(N__11152),
            .in2(_gnd_net_),
            .in3(N__11032),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_2 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_1 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_2 ),
            .clk(N__29453),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_3_LC_1_6_2 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_3_LC_1_6_2 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_3_LC_1_6_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_3_LC_1_6_2  (
            .in0(N__11524),
            .in1(N__11161),
            .in2(_gnd_net_),
            .in3(N__11212),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_3 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_2 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_3 ),
            .clk(N__29453),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_4_LC_1_6_3 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_4_LC_1_6_3 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_4_LC_1_6_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_4_LC_1_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11188),
            .in3(N__11209),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_4 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_3 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_4 ),
            .clk(N__29453),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_5_LC_1_6_4 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_5_LC_1_6_4 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_5_LC_1_6_4 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_5_LC_1_6_4  (
            .in0(N__11525),
            .in1(_gnd_net_),
            .in2(N__11200),
            .in3(N__11206),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_5 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_4 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_5 ),
            .clk(N__29453),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_6_LC_1_6_5 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_6_LC_1_6_5 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_6_LC_1_6_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_6_LC_1_6_5  (
            .in0(N__11175),
            .in1(N__11523),
            .in2(_gnd_net_),
            .in3(N__11203),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29453),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_RNII048_6_LC_1_6_6 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_RNII048_6_LC_1_6_6 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.counter_RNII048_6_LC_1_6_6 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_RNII048_6_LC_1_6_6  (
            .in0(N__11196),
            .in1(N__11184),
            .in2(N__11176),
            .in3(N__11160),
            .lcout(),
            .ltout(\buart.Z_tx.Z_baudgen.ser_clk_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_1_6_7 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_1_6_7 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_1_6_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_1_6_7  (
            .in0(N__11119),
            .in1(N__11151),
            .in2(N__11143),
            .in3(N__11135),
            .lcout(\buart.Z_tx.ser_clk ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_1_LC_1_7_2 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_1_LC_1_7_2 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_1_LC_1_7_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_1_LC_1_7_2  (
            .in0(N__11122),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11139),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29445),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_0_LC_1_7_5 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_0_LC_1_7_5 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_0_LC_1_7_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_0_LC_1_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11121),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29445),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_0_ret_29_RNO_2_LC_1_10_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_29_RNO_2_LC_1_10_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_0_ret_29_RNO_2_LC_1_10_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_29_RNO_2_LC_1_10_0  (
            .in0(N__21576),
            .in1(N__15472),
            .in2(N__17565),
            .in3(N__15377),
            .lcout(\Lab_UT.dictrl.N_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_0_ret_29_RNO_4_LC_1_10_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_29_RNO_4_LC_1_10_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_0_ret_29_RNO_4_LC_1_10_1 .LUT_INIT=16'b0001011100000000;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_29_RNO_4_LC_1_10_1  (
            .in0(N__20813),
            .in1(N__21577),
            .in2(N__11236),
            .in3(N__21110),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_17_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_0_ret_29_RNO_1_LC_1_10_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_29_RNO_1_LC_1_10_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_0_ret_29_RNO_1_LC_1_10_2 .LUT_INIT=16'b1111111011110000;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_29_RNO_1_LC_1_10_2  (
            .in0(N__21111),
            .in1(N__15473),
            .in2(N__11248),
            .in3(N__11224),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_i_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_0_ret_29_LC_1_10_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_29_LC_1_10_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.currState_0_ret_29_LC_1_10_3 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_29_LC_1_10_3  (
            .in0(N__17137),
            .in1(N__24681),
            .in2(N__11245),
            .in3(N__11242),
            .lcout(Lab_UT_dictrl_r_Sone_init17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29422),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_RNIN0MBN_1_LC_1_10_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_RNIN0MBN_1_LC_1_10_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_RNIN0MBN_1_LC_1_10_4 .LUT_INIT=16'b0011011100110010;
    LogicCell40 \Lab_UT.dictrl.currState_2_RNIN0MBN_1_LC_1_10_4  (
            .in0(N__23345),
            .in1(N__11218),
            .in2(N__17929),
            .in3(N__17231),
            .lcout(\Lab_UT.dictrl.N_8_2 ),
            .ltout(\Lab_UT.dictrl.N_8_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_0_ret_29_RNO_3_LC_1_10_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_29_RNO_3_LC_1_10_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_0_ret_29_RNO_3_LC_1_10_5 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_29_RNO_3_LC_1_10_5  (
            .in0(_gnd_net_),
            .in1(N__17548),
            .in2(N__11227),
            .in3(N__21575),
            .lcout(\Lab_UT.dictrl.g0_i_a8_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_RNIGHD18_0_1_LC_1_10_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_RNIGHD18_0_1_LC_1_10_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_RNIGHD18_0_1_LC_1_10_6 .LUT_INIT=16'b0101010111110000;
    LogicCell40 \Lab_UT.dictrl.nextState_RNIGHD18_0_1_LC_1_10_6  (
            .in0(N__13863),
            .in1(_gnd_net_),
            .in2(N__13834),
            .in3(N__18063),
            .lcout(\Lab_UT.dictrl.N_1605_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_RNO_12_1_LC_1_10_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_RNO_12_1_LC_1_10_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_RNO_12_1_LC_1_10_7 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \Lab_UT.dictrl.nextState_RNO_12_1_LC_1_10_7  (
            .in0(N__18064),
            .in1(N__13830),
            .in2(_gnd_net_),
            .in3(N__13862),
            .lcout(\Lab_UT.dictrl.N_1605_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_RNO_7_1_LC_1_11_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_RNO_7_1_LC_1_11_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_RNO_7_1_LC_1_11_0 .LUT_INIT=16'b0011011100110010;
    LogicCell40 \Lab_UT.dictrl.nextState_RNO_7_1_LC_1_11_0  (
            .in0(N__23376),
            .in1(N__17304),
            .in2(N__17893),
            .in3(N__17258),
            .lcout(\Lab_UT.dictrl.N_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_0_ret_0_LC_1_11_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_0_LC_1_11_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.currState_0_ret_0_LC_1_11_1 .LUT_INIT=16'b1110110011101111;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_0_LC_1_11_1  (
            .in0(N__17260),
            .in1(N__24671),
            .in2(N__17181),
            .in3(N__17303),
            .lcout(\Lab_UT.dictrl.currState_i_5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29413),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_0_ret_28_RNO_4_LC_1_11_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_28_RNO_4_LC_1_11_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_0_ret_28_RNO_4_LC_1_11_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_28_RNO_4_LC_1_11_2  (
            .in0(_gnd_net_),
            .in1(N__23375),
            .in2(_gnd_net_),
            .in3(N__17828),
            .lcout(),
            .ltout(\Lab_UT.dictrl.currState_0_ret_28_RNOZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_0_ret_28_RNO_2_LC_1_11_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_28_RNO_2_LC_1_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_0_ret_28_RNO_2_LC_1_11_3 .LUT_INIT=16'b1111111110100011;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_28_RNO_2_LC_1_11_3  (
            .in0(N__17259),
            .in1(N__17302),
            .in2(N__11299),
            .in3(N__24669),
            .lcout(\Lab_UT.dictrl.currState_0_ret_28_RNOZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_RNO_6_1_LC_1_11_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_RNO_6_1_LC_1_11_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_RNO_6_1_LC_1_11_4 .LUT_INIT=16'b0011011100110010;
    LogicCell40 \Lab_UT.dictrl.nextState_RNO_6_1_LC_1_11_4  (
            .in0(N__23377),
            .in1(N__11296),
            .in2(N__17894),
            .in3(N__17257),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_RNO_2_1_LC_1_11_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_RNO_2_1_LC_1_11_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_RNO_2_1_LC_1_11_5 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \Lab_UT.dictrl.nextState_RNO_2_1_LC_1_11_5  (
            .in0(N__11290),
            .in1(N__15476),
            .in2(N__11284),
            .in3(N__21112),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_i_o4_4_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_RNO_0_1_LC_1_11_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_RNO_0_1_LC_1_11_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_RNO_0_1_LC_1_11_6 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \Lab_UT.dictrl.nextState_RNO_0_1_LC_1_11_6  (
            .in0(N__24670),
            .in1(N__17572),
            .in2(N__11281),
            .in3(N__21625),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_i_o4_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_LC_1_11_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_LC_1_11_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.nextState_1_LC_1_11_7 .LUT_INIT=16'b1010101010100011;
    LogicCell40 \Lab_UT.dictrl.nextState_1_LC_1_11_7  (
            .in0(N__13223),
            .in1(N__12277),
            .in2(N__11278),
            .in3(N__15253),
            .lcout(\Lab_UT.dictrl.nextState_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29413),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.hh_0_LC_1_12_3 .C_ON=1'b0;
    defparam \buart.Z_rx.hh_0_LC_1_12_3 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.hh_0_LC_1_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.hh_0_LC_1_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11275),
            .lcout(\buart.Z_rx.hhZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29405),
            .ce(),
            .sr(N__26078));
    defparam \uu0.l_count_RNI04591_10_LC_2_1_0 .C_ON=1'b0;
    defparam \uu0.l_count_RNI04591_10_LC_2_1_0 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNI04591_10_LC_2_1_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uu0.l_count_RNI04591_10_LC_2_1_0  (
            .in0(N__11266),
            .in1(N__11321),
            .in2(N__11347),
            .in3(N__11395),
            .lcout(),
            .ltout(\uu0.un4_l_count_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_RNI2GS72_4_LC_2_1_1 .C_ON=1'b0;
    defparam \uu0.l_count_RNI2GS72_4_LC_2_1_1 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNI2GS72_4_LC_2_1_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \uu0.l_count_RNI2GS72_4_LC_2_1_1  (
            .in0(N__12513),
            .in1(N__12474),
            .in2(N__11251),
            .in3(N__11360),
            .lcout(),
            .ltout(\uu0.un4_l_count_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_RNI8ORT6_11_LC_2_1_2 .C_ON=1'b0;
    defparam \uu0.l_count_RNI8ORT6_11_LC_2_1_2 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNI8ORT6_11_LC_2_1_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.l_count_RNI8ORT6_11_LC_2_1_2  (
            .in0(N__11437),
            .in1(N__11575),
            .in2(N__11431),
            .in3(N__11782),
            .lcout(\uu0.un4_l_count_0 ),
            .ltout(\uu0.un4_l_count_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_11_LC_2_1_3 .C_ON=1'b0;
    defparam \uu0.l_count_11_LC_2_1_3 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_11_LC_2_1_3 .LUT_INIT=16'b0000011100001000;
    LogicCell40 \uu0.l_count_11_LC_2_1_3  (
            .in0(N__11723),
            .in1(N__11425),
            .in2(N__11428),
            .in3(N__11418),
            .lcout(\uu0.l_countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29479),
            .ce(N__12345),
            .sr(N__26088));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_2_1_4 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_2_1_4 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_2_1_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_2_1_4  (
            .in0(N__11640),
            .in1(N__11323),
            .in2(_gnd_net_),
            .in3(N__11397),
            .lcout(\uu0.un143_ci_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_10_LC_2_1_5 .C_ON=1'b0;
    defparam \uu0.l_count_10_LC_2_1_5 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_10_LC_2_1_5 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu0.l_count_10_LC_2_1_5  (
            .in0(N__11725),
            .in1(N__11641),
            .in2(N__11401),
            .in3(N__11326),
            .lcout(\uu0.l_countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29479),
            .ce(N__12345),
            .sr(N__26088));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_2_1_6 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_2_1_6 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_2_1_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_2_1_6  (
            .in0(N__11639),
            .in1(N__11322),
            .in2(N__11419),
            .in3(N__11396),
            .lcout(\uu0.un154_ci_9 ),
            .ltout(\uu0.un154_ci_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_14_LC_2_1_7 .C_ON=1'b0;
    defparam \uu0.l_count_14_LC_2_1_7 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_14_LC_2_1_7 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu0.l_count_14_LC_2_1_7  (
            .in0(N__11724),
            .in1(N__11344),
            .in2(N__11365),
            .in3(N__11361),
            .lcout(\uu0.l_countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29479),
            .ce(N__12345),
            .sr(N__26088));
    defparam \uu0.l_count_9_LC_2_2_0 .C_ON=1'b0;
    defparam \uu0.l_count_9_LC_2_2_0 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_9_LC_2_2_0 .LUT_INIT=16'b0011111111000000;
    LogicCell40 \uu0.l_count_9_LC_2_2_0  (
            .in0(_gnd_net_),
            .in1(N__11324),
            .in2(N__11735),
            .in3(N__11638),
            .lcout(\uu0.l_countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29475),
            .ce(N__12344),
            .sr(N__26086));
    defparam \uu0.l_count_8_LC_2_2_1 .C_ON=1'b0;
    defparam \uu0.l_count_8_LC_2_2_1 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_8_LC_2_2_1 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \uu0.l_count_8_LC_2_2_1  (
            .in0(N__11325),
            .in1(N__11716),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uu0.l_countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29475),
            .ce(N__12344),
            .sr(N__26086));
    defparam \uu0.l_count_17_LC_2_2_2 .C_ON=1'b0;
    defparam \uu0.l_count_17_LC_2_2_2 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_17_LC_2_2_2 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu0.l_count_17_LC_2_2_2  (
            .in0(N__11683),
            .in1(N__11604),
            .in2(N__11734),
            .in3(N__11662),
            .lcout(\uu0.l_countZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29475),
            .ce(N__12344),
            .sr(N__26086));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_2_2_3 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_2_2_3 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_2_2_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_2_2_3  (
            .in0(N__12400),
            .in1(N__12379),
            .in2(N__12433),
            .in3(N__11616),
            .lcout(\uu0.un110_ci ),
            .ltout(\uu0.un110_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_2_2_4 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_2_2_4 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_2_2_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_2_2_4  (
            .in0(N__11682),
            .in1(N__11603),
            .in2(N__11665),
            .in3(N__11661),
            .lcout(),
            .ltout(\uu0.un220_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_18_LC_2_2_5 .C_ON=1'b0;
    defparam \uu0.l_count_18_LC_2_2_5 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_18_LC_2_2_5 .LUT_INIT=16'b0000000000111100;
    LogicCell40 \uu0.l_count_18_LC_2_2_5  (
            .in0(_gnd_net_),
            .in1(N__11815),
            .in2(N__11644),
            .in3(N__12985),
            .lcout(\uu0.l_countZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29475),
            .ce(N__12344),
            .sr(N__26086));
    defparam \uu0.l_count_7_LC_2_2_6 .C_ON=1'b0;
    defparam \uu0.l_count_7_LC_2_2_6 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_7_LC_2_2_6 .LUT_INIT=16'b0001010001010000;
    LogicCell40 \uu0.l_count_7_LC_2_2_6  (
            .in0(N__12986),
            .in1(N__12493),
            .in2(N__11620),
            .in3(N__12401),
            .lcout(\uu0.l_countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29475),
            .ce(N__12344),
            .sr(N__26086));
    defparam \uu0.l_count_RNIRLTJ1_17_LC_2_2_7 .C_ON=1'b0;
    defparam \uu0.l_count_RNIRLTJ1_17_LC_2_2_7 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNIRLTJ1_17_LC_2_2_7 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \uu0.l_count_RNIRLTJ1_17_LC_2_2_7  (
            .in0(N__11637),
            .in1(N__11615),
            .in2(N__11605),
            .in3(N__11588),
            .lcout(\uu0.un4_l_count_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_0_LC_2_3_1 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_0_LC_2_3_1 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.bitcount_0_LC_2_3_1 .LUT_INIT=16'b0000011000001010;
    LogicCell40 \buart.Z_tx.bitcount_0_LC_2_3_1  (
            .in0(N__11480),
            .in1(N__11569),
            .in2(N__12832),
            .in3(N__11530),
            .lcout(\buart.Z_tx.bitcountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29469),
            .ce(),
            .sr(N__26084));
    defparam \uu0.delay_line_0_LC_2_3_2 .C_ON=1'b0;
    defparam \uu0.delay_line_0_LC_2_3_2 .SEQ_MODE=4'b1010;
    defparam \uu0.delay_line_0_LC_2_3_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.delay_line_0_LC_2_3_2  (
            .in0(N__11869),
            .in1(N__12523),
            .in2(N__11854),
            .in3(N__11455),
            .lcout(\uu0.delay_lineZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29469),
            .ce(),
            .sr(N__26084));
    defparam \uu0.l_precount_3_LC_2_3_3 .C_ON=1'b0;
    defparam \uu0.l_precount_3_LC_2_3_3 .SEQ_MODE=4'b1010;
    defparam \uu0.l_precount_3_LC_2_3_3 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu0.l_precount_3_LC_2_3_3  (
            .in0(N__11457),
            .in1(N__11852),
            .in2(N__12529),
            .in3(N__11872),
            .lcout(\uu0.l_precountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29469),
            .ce(),
            .sr(N__26084));
    defparam \uu0.l_precount_2_LC_2_3_4 .C_ON=1'b0;
    defparam \uu0.l_precount_2_LC_2_3_4 .SEQ_MODE=4'b1010;
    defparam \uu0.l_precount_2_LC_2_3_4 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \uu0.l_precount_2_LC_2_3_4  (
            .in0(N__11871),
            .in1(N__12525),
            .in2(_gnd_net_),
            .in3(N__11456),
            .lcout(\uu0.l_precountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29469),
            .ce(),
            .sr(N__26084));
    defparam \uu0.l_precount_1_LC_2_3_5 .C_ON=1'b0;
    defparam \uu0.l_precount_1_LC_2_3_5 .SEQ_MODE=4'b1010;
    defparam \uu0.l_precount_1_LC_2_3_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \uu0.l_precount_1_LC_2_3_5  (
            .in0(N__12524),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11870),
            .lcout(\uu0.l_precountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29469),
            .ce(),
            .sr(N__26084));
    defparam \uu0.l_precount_RNI85Q91_3_LC_2_3_6 .C_ON=1'b0;
    defparam \uu0.l_precount_RNI85Q91_3_LC_2_3_6 .SEQ_MODE=4'b0000;
    defparam \uu0.l_precount_RNI85Q91_3_LC_2_3_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uu0.l_precount_RNI85Q91_3_LC_2_3_6  (
            .in0(N__11868),
            .in1(N__12451),
            .in2(N__11853),
            .in3(N__11830),
            .lcout(),
            .ltout(\uu0.un4_l_count_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_RNI96A32_18_LC_2_3_7 .C_ON=1'b0;
    defparam \uu0.l_count_RNI96A32_18_LC_2_3_7 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNI96A32_18_LC_2_3_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.l_count_RNI96A32_18_LC_2_3_7  (
            .in0(N__11814),
            .in1(N__11803),
            .in2(N__11785),
            .in3(N__12375),
            .lcout(\uu0.un4_l_count_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_0_LC_2_4_0 .C_ON=1'b0;
    defparam \uu2.r_data_reg_0_LC_2_4_0 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_0_LC_2_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_0_LC_2_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11773),
            .lcout(vbuf_tx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__12595),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_1_LC_2_4_1 .C_ON=1'b0;
    defparam \uu2.r_data_reg_1_LC_2_4_1 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_1_LC_2_4_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_1_LC_2_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11767),
            .lcout(vbuf_tx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__12595),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_2_LC_2_4_2 .C_ON=1'b0;
    defparam \uu2.r_data_reg_2_LC_2_4_2 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_2_LC_2_4_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_2_LC_2_4_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11761),
            .lcout(vbuf_tx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__12595),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_3_LC_2_4_3 .C_ON=1'b0;
    defparam \uu2.r_data_reg_3_LC_2_4_3 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_3_LC_2_4_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_3_LC_2_4_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11755),
            .lcout(vbuf_tx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__12595),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_4_LC_2_4_4 .C_ON=1'b0;
    defparam \uu2.r_data_reg_4_LC_2_4_4 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_4_LC_2_4_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_4_LC_2_4_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11749),
            .lcout(vbuf_tx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__12595),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_5_LC_2_4_5 .C_ON=1'b0;
    defparam \uu2.r_data_reg_5_LC_2_4_5 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_5_LC_2_4_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uu2.r_data_reg_5_LC_2_4_5  (
            .in0(N__11743),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(vbuf_tx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__12595),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_6_LC_2_4_6 .C_ON=1'b0;
    defparam \uu2.r_data_reg_6_LC_2_4_6 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_6_LC_2_4_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_6_LC_2_4_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11953),
            .lcout(vbuf_tx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__12595),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_7_LC_2_4_7 .C_ON=1'b0;
    defparam \uu2.r_data_reg_7_LC_2_4_7 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_7_LC_2_4_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_7_LC_2_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11947),
            .lcout(vbuf_tx_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__12595),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_1_LC_2_5_0 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_1_LC_2_5_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_1_LC_2_5_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \buart.Z_tx.shifter_1_LC_2_5_0  (
            .in0(N__11941),
            .in1(N__11902),
            .in2(_gnd_net_),
            .in3(N__12816),
            .lcout(\buart.Z_tx.shifterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29454),
            .ce(N__12729),
            .sr(N__26080));
    defparam \buart.Z_tx.shifter_0_LC_2_5_1 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_0_LC_2_5_1 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_0_LC_2_5_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \buart.Z_tx.shifter_0_LC_2_5_1  (
            .in0(N__12812),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11935),
            .lcout(\buart.Z_tx.shifterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29454),
            .ce(N__12729),
            .sr(N__26080));
    defparam \buart.Z_tx.uart_tx_LC_2_5_2 .C_ON=1'b0;
    defparam \buart.Z_tx.uart_tx_LC_2_5_2 .SEQ_MODE=4'b1011;
    defparam \buart.Z_tx.uart_tx_LC_2_5_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \buart.Z_tx.uart_tx_LC_2_5_2  (
            .in0(_gnd_net_),
            .in1(N__11929),
            .in2(_gnd_net_),
            .in3(N__12819),
            .lcout(o_serial_data_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29454),
            .ce(N__12729),
            .sr(N__26080));
    defparam \buart.Z_tx.shifter_2_LC_2_5_3 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_2_LC_2_5_3 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_2_LC_2_5_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \buart.Z_tx.shifter_2_LC_2_5_3  (
            .in0(N__12813),
            .in1(N__11890),
            .in2(_gnd_net_),
            .in3(N__11908),
            .lcout(\buart.Z_tx.shifterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29454),
            .ce(N__12729),
            .sr(N__26080));
    defparam \buart.Z_tx.shifter_3_LC_2_5_4 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_3_LC_2_5_4 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_3_LC_2_5_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \buart.Z_tx.shifter_3_LC_2_5_4  (
            .in0(N__11878),
            .in1(N__12817),
            .in2(_gnd_net_),
            .in3(N__11896),
            .lcout(\buart.Z_tx.shifterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29454),
            .ce(N__12729),
            .sr(N__26080));
    defparam \buart.Z_tx.shifter_4_LC_2_5_5 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_4_LC_2_5_5 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_4_LC_2_5_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \buart.Z_tx.shifter_4_LC_2_5_5  (
            .in0(N__12814),
            .in1(N__11986),
            .in2(_gnd_net_),
            .in3(N__11884),
            .lcout(\buart.Z_tx.shifterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29454),
            .ce(N__12729),
            .sr(N__26080));
    defparam \buart.Z_tx.shifter_5_LC_2_5_6 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_5_LC_2_5_6 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_5_LC_2_5_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \buart.Z_tx.shifter_5_LC_2_5_6  (
            .in0(N__11974),
            .in1(N__12818),
            .in2(_gnd_net_),
            .in3(N__11992),
            .lcout(\buart.Z_tx.shifterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29454),
            .ce(N__12729),
            .sr(N__26080));
    defparam \buart.Z_tx.shifter_6_LC_2_5_7 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_6_LC_2_5_7 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_6_LC_2_5_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \buart.Z_tx.shifter_6_LC_2_5_7  (
            .in0(N__12815),
            .in1(N__12844),
            .in2(_gnd_net_),
            .in3(N__11980),
            .lcout(\buart.Z_tx.shifterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29454),
            .ce(N__12729),
            .sr(N__26080));
    defparam \uu2.vram_rd_clk_det_0_LC_2_6_0 .C_ON=1'b0;
    defparam \uu2.vram_rd_clk_det_0_LC_2_6_0 .SEQ_MODE=4'b1011;
    defparam \uu2.vram_rd_clk_det_0_LC_2_6_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.vram_rd_clk_det_0_LC_2_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13466),
            .lcout(\uu2.vram_rd_clk_detZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.vram_rd_clk_det_0C_net ),
            .ce(),
            .sr(N__26050));
    defparam \uu2.vram_rd_clk_det_1_LC_2_6_1 .C_ON=1'b0;
    defparam \uu2.vram_rd_clk_det_1_LC_2_6_1 .SEQ_MODE=4'b1011;
    defparam \uu2.vram_rd_clk_det_1_LC_2_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.vram_rd_clk_det_1_LC_2_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12609),
            .lcout(\uu2.vram_rd_clk_detZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.vram_rd_clk_det_0C_net ),
            .ce(),
            .sr(N__26050));
    defparam \uu2.l_count_3_LC_2_7_0 .C_ON=1'b0;
    defparam \uu2.l_count_3_LC_2_7_0 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_3_LC_2_7_0 .LUT_INIT=16'b0001001100100000;
    LogicCell40 \uu2.l_count_3_LC_2_7_0  (
            .in0(N__12127),
            .in1(N__12938),
            .in2(N__13048),
            .in3(N__12109),
            .lcout(\uu2.l_countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29438),
            .ce(),
            .sr(N__26077));
    defparam \uu2.l_count_2_LC_2_7_1 .C_ON=1'b0;
    defparam \uu2.l_count_2_LC_2_7_1 .SEQ_MODE=4'b1011;
    defparam \uu2.l_count_2_LC_2_7_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.l_count_2_LC_2_7_1  (
            .in0(_gnd_net_),
            .in1(N__13044),
            .in2(_gnd_net_),
            .in3(N__12126),
            .lcout(\uu2.l_countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29438),
            .ce(),
            .sr(N__26077));
    defparam \uu2.l_count_RNIFGGK1_3_LC_2_7_2 .C_ON=1'b0;
    defparam \uu2.l_count_RNIFGGK1_3_LC_2_7_2 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNIFGGK1_3_LC_2_7_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uu2.l_count_RNIFGGK1_3_LC_2_7_2  (
            .in0(N__12005),
            .in1(N__12056),
            .in2(N__12079),
            .in3(N__12107),
            .lcout(\uu2.un1_l_count_1_3 ),
            .ltout(\uu2.un1_l_count_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_RNI9S834_0_1_LC_2_7_3 .C_ON=1'b0;
    defparam \uu2.l_count_RNI9S834_0_1_LC_2_7_3 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNI9S834_0_1_LC_2_7_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.l_count_RNI9S834_0_1_LC_2_7_3  (
            .in0(N__13116),
            .in1(N__12124),
            .in2(N__11968),
            .in3(N__12091),
            .lcout(\uu2.un1_l_count_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_RNI9S834_1_LC_2_7_4 .C_ON=1'b0;
    defparam \uu2.l_count_RNI9S834_1_LC_2_7_4 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNI9S834_1_LC_2_7_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.l_count_RNI9S834_1_LC_2_7_4  (
            .in0(N__12125),
            .in1(N__12145),
            .in2(N__11965),
            .in3(N__13117),
            .lcout(\uu2.un1_l_count_2_0 ),
            .ltout(\uu2.un1_l_count_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_4_LC_2_7_5 .C_ON=1'b0;
    defparam \uu2.l_count_4_LC_2_7_5 .SEQ_MODE=4'b1011;
    defparam \uu2.l_count_4_LC_2_7_5 .LUT_INIT=16'b0000001100001100;
    LogicCell40 \uu2.l_count_4_LC_2_7_5  (
            .in0(_gnd_net_),
            .in1(N__12025),
            .in2(N__11956),
            .in3(N__12182),
            .lcout(\uu2.l_countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29438),
            .ce(),
            .sr(N__26077));
    defparam \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_2_7_6 .C_ON=1'b0;
    defparam \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_2_7_6 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_2_7_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_2_7_6  (
            .in0(N__12123),
            .in1(N__12108),
            .in2(N__13090),
            .in3(N__13115),
            .lcout(\uu2.un306_ci ),
            .ltout(\uu2.un306_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_5_LC_2_7_7 .C_ON=1'b0;
    defparam \uu2.l_count_5_LC_2_7_7 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_5_LC_2_7_7 .LUT_INIT=16'b0101101010101010;
    LogicCell40 \uu2.l_count_5_LC_2_7_7  (
            .in0(N__12057),
            .in1(_gnd_net_),
            .in2(N__12097),
            .in3(N__12183),
            .lcout(\uu2.l_countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29438),
            .ce(),
            .sr(N__26077));
    defparam \uu2.vbuf_count.counter_gen_label_8__un350_ci_LC_2_8_0 .C_ON=1'b0;
    defparam \uu2.vbuf_count.counter_gen_label_8__un350_ci_LC_2_8_0 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_count.counter_gen_label_8__un350_ci_LC_2_8_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.vbuf_count.counter_gen_label_8__un350_ci_LC_2_8_0  (
            .in0(N__12200),
            .in1(N__12006),
            .in2(N__12042),
            .in3(N__12022),
            .lcout(\uu2.un350_ci ),
            .ltout(\uu2.un350_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_9_LC_2_8_1 .C_ON=1'b0;
    defparam \uu2.l_count_9_LC_2_8_1 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_9_LC_2_8_1 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \uu2.l_count_9_LC_2_8_1  (
            .in0(N__12078),
            .in1(N__12159),
            .in2(N__12094),
            .in3(N__12939),
            .lcout(\uu2.l_countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29431),
            .ce(),
            .sr(N__26076));
    defparam \uu2.l_count_RNIBCGK1_0_9_LC_2_8_2 .C_ON=1'b0;
    defparam \uu2.l_count_RNIBCGK1_0_9_LC_2_8_2 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNIBCGK1_0_9_LC_2_8_2 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \uu2.l_count_RNIBCGK1_0_9_LC_2_8_2  (
            .in0(N__12198),
            .in1(N__12177),
            .in2(N__12160),
            .in3(N__13088),
            .lcout(\uu2.un1_l_count_1_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_8_LC_2_8_3 .C_ON=1'b0;
    defparam \uu2.l_count_8_LC_2_8_3 .SEQ_MODE=4'b1011;
    defparam \uu2.l_count_8_LC_2_8_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.l_count_8_LC_2_8_3  (
            .in0(_gnd_net_),
            .in1(N__12077),
            .in2(_gnd_net_),
            .in3(N__12085),
            .lcout(\uu2.l_countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29431),
            .ce(),
            .sr(N__26076));
    defparam \uu2.l_count_6_LC_2_8_4 .C_ON=1'b0;
    defparam \uu2.l_count_6_LC_2_8_4 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_6_LC_2_8_4 .LUT_INIT=16'b0101101010101010;
    LogicCell40 \uu2.l_count_6_LC_2_8_4  (
            .in0(N__12201),
            .in1(_gnd_net_),
            .in2(N__12043),
            .in3(N__12023),
            .lcout(\uu2.l_countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29431),
            .ce(),
            .sr(N__26076));
    defparam \uu2.vbuf_count.counter_gen_label_6__un328_ci_3_LC_2_8_5 .C_ON=1'b0;
    defparam \uu2.vbuf_count.counter_gen_label_6__un328_ci_3_LC_2_8_5 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_count.counter_gen_label_6__un328_ci_3_LC_2_8_5 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \uu2.vbuf_count.counter_gen_label_6__un328_ci_3_LC_2_8_5  (
            .in0(N__12181),
            .in1(N__12058),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uu2.vbuf_count.un328_ci_3 ),
            .ltout(\uu2.vbuf_count.un328_ci_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_7_LC_2_8_6 .C_ON=1'b0;
    defparam \uu2.l_count_7_LC_2_8_6 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_7_LC_2_8_6 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu2.l_count_7_LC_2_8_6  (
            .in0(N__12202),
            .in1(N__12007),
            .in2(N__12028),
            .in3(N__12024),
            .lcout(\uu2.l_countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29431),
            .ce(),
            .sr(N__26076));
    defparam \uu2.l_count_RNIBCGK1_9_LC_2_8_7 .C_ON=1'b0;
    defparam \uu2.l_count_RNIBCGK1_9_LC_2_8_7 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNIBCGK1_9_LC_2_8_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \uu2.l_count_RNIBCGK1_9_LC_2_8_7  (
            .in0(N__13089),
            .in1(N__12199),
            .in2(N__12184),
            .in3(N__12158),
            .lcout(\uu2.un1_l_count_2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_0_rep2_RNIOBFP3_LC_2_9_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_0_rep2_RNIOBFP3_LC_2_9_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_0_rep2_RNIOBFP3_LC_2_9_0 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \Lab_UT.dictrl.currState_2_0_rep2_RNIOBFP3_LC_2_9_0  (
            .in0(N__24878),
            .in1(N__27790),
            .in2(N__20950),
            .in3(N__27542),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_8_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_RNIA5707_2_LC_2_9_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_RNIA5707_2_LC_2_9_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_RNIA5707_2_LC_2_9_1 .LUT_INIT=16'b0100000011001000;
    LogicCell40 \Lab_UT.dictrl.currState_2_RNIA5707_2_LC_2_9_1  (
            .in0(N__25020),
            .in1(N__12214),
            .in2(N__12139),
            .in3(N__12133),
            .lcout(\Lab_UT.dictrl.N_23_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_13_LC_2_9_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_13_LC_2_9_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_13_LC_2_9_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__g0_13_LC_2_9_2  (
            .in0(N__20949),
            .in1(N__27789),
            .in2(_gnd_net_),
            .in3(N__27541),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_20_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_5_LC_2_9_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_5_LC_2_9_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_5_LC_2_9_3 .LUT_INIT=16'b0100011111001111;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__g0_5_LC_2_9_3  (
            .in0(N__21245),
            .in1(N__23826),
            .in2(N__12136),
            .in3(N__17112),
            .lcout(\Lab_UT.dictrl.N_30_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_RNIKTU5_2_LC_2_9_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_RNIKTU5_2_LC_2_9_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_RNIKTU5_2_LC_2_9_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.dictrl.nextState_RNIKTU5_2_LC_2_9_4  (
            .in0(_gnd_net_),
            .in1(N__15541),
            .in2(_gnd_net_),
            .in3(N__23326),
            .lcout(\Lab_UT.dictrl.G_19_0_a7_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_0_ret_21_RNI40BJ2_LC_2_9_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_21_RNI40BJ2_LC_2_9_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_0_ret_21_RNI40BJ2_LC_2_9_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_21_RNI40BJ2_LC_2_9_5  (
            .in0(N__27296),
            .in1(N__20361),
            .in2(_gnd_net_),
            .in3(N__24005),
            .lcout(\Lab_UT.dictrl.N_9_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_3_3_rep1_RNIO9JG3_LC_2_9_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_3_3_rep1_RNIO9JG3_LC_2_9_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_3_3_rep1_RNIO9JG3_LC_2_9_6 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \Lab_UT.dictrl.currState_3_3_rep1_RNIO9JG3_LC_2_9_6  (
            .in0(N__20360),
            .in1(N__27297),
            .in2(N__14269),
            .in3(N__23327),
            .lcout(\Lab_UT.dictrl.G_30_0_a7_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_fast_RNI13TV_0_LC_2_9_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_fast_RNI13TV_0_LC_2_9_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_fast_RNI13TV_0_LC_2_9_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \Lab_UT.dictrl.currState_2_fast_RNI13TV_0_LC_2_9_7  (
            .in0(N__25019),
            .in1(N__17861),
            .in2(N__24897),
            .in3(N__14500),
            .lcout(\Lab_UT.dictrl.G_30_0_a7_4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_0_ret_29_RNIK6A94_LC_2_10_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_29_RNIK6A94_LC_2_10_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_0_ret_29_RNIK6A94_LC_2_10_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_29_RNIK6A94_LC_2_10_0  (
            .in0(N__27561),
            .in1(N__27809),
            .in2(N__12253),
            .in3(N__23341),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_31_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_0_ret_29_RNINPDOC_LC_2_10_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_29_RNINPDOC_LC_2_10_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_0_ret_29_RNINPDOC_LC_2_10_1 .LUT_INIT=16'b1111111111110010;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_29_RNINPDOC_LC_2_10_1  (
            .in0(N__12244),
            .in1(N__12271),
            .in2(N__12238),
            .in3(N__12220),
            .lcout(),
            .ltout(\Lab_UT.dictrl.G_30_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_0_ret_21_RNI66NNS_LC_2_10_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_21_RNI66NNS_LC_2_10_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_0_ret_21_RNI66NNS_LC_2_10_2 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_21_RNI66NNS_LC_2_10_2  (
            .in0(N__12265),
            .in1(N__12235),
            .in2(N__12229),
            .in3(N__21133),
            .lcout(\Lab_UT.dictrl.nextStateZ0Z_1 ),
            .ltout(\Lab_UT.dictrl.nextStateZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_0_ret_21_RNIAVHPS_LC_2_10_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_21_RNIAVHPS_LC_2_10_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_0_ret_21_RNIAVHPS_LC_2_10_3 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_21_RNIAVHPS_LC_2_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12226),
            .in3(N__24680),
            .lcout(\Lab_UT.dictrl.N_10ctr ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_3_3_rep1_RNIPTVF_LC_2_10_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_3_3_rep1_RNIPTVF_LC_2_10_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_3_3_rep1_RNIPTVF_LC_2_10_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Lab_UT.dictrl.currState_3_3_rep1_RNIPTVF_LC_2_10_4  (
            .in0(_gnd_net_),
            .in1(N__17860),
            .in2(_gnd_net_),
            .in3(N__20334),
            .lcout(),
            .ltout(\Lab_UT.dictrl.G_30_0_a7_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_RNIO37J1_1_LC_2_10_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_RNIO37J1_1_LC_2_10_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_RNIO37J1_1_LC_2_10_5 .LUT_INIT=16'b1101100010001000;
    LogicCell40 \Lab_UT.dictrl.nextState_RNIO37J1_1_LC_2_10_5  (
            .in0(N__23343),
            .in1(N__13216),
            .in2(N__12223),
            .in3(N__14268),
            .lcout(\Lab_UT.dictrl.G_30_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_RNI1O2A_1_LC_2_10_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_RNI1O2A_1_LC_2_10_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_RNI1O2A_1_LC_2_10_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Lab_UT.dictrl.currState_2_RNI1O2A_1_LC_2_10_6  (
            .in0(_gnd_net_),
            .in1(N__17859),
            .in2(_gnd_net_),
            .in3(N__23340),
            .lcout(\Lab_UT.dictrl.G_30_0_a7_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_RNI0P25D_1_LC_2_10_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_RNI0P25D_1_LC_2_10_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_RNI0P25D_1_LC_2_10_7 .LUT_INIT=16'b1011000011110100;
    LogicCell40 \Lab_UT.dictrl.currState_2_RNI0P25D_1_LC_2_10_7  (
            .in0(N__23342),
            .in1(N__17862),
            .in2(N__15157),
            .in3(N__12208),
            .lcout(\Lab_UT.dictrl.currState_2_RNI0P25DZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_0_LC_2_11_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_0_LC_2_11_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_0_LC_2_11_0 .LUT_INIT=16'b1101100010001000;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__g0_0_LC_2_11_0  (
            .in0(N__25045),
            .in1(N__13864),
            .in2(N__24899),
            .in3(N__15336),
            .lcout(),
            .ltout(\Lab_UT.dictrl.i8_mux_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_LC_2_11_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_LC_2_11_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_LC_2_11_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__g0_LC_2_11_1  (
            .in0(N__17888),
            .in1(_gnd_net_),
            .in2(N__12280),
            .in3(N__17261),
            .lcout(\Lab_UT.dictrl.i7_mux_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_RNIJ59B3_2_LC_2_11_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_RNIJ59B3_2_LC_2_11_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_RNIJ59B3_2_LC_2_11_2 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \Lab_UT.dictrl.currState_2_RNIJ59B3_2_LC_2_11_2  (
            .in0(N__25041),
            .in1(N__17886),
            .in2(N__24898),
            .in3(N__27543),
            .lcout(\Lab_UT.dictrl.N_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_1_LC_2_11_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_1_LC_2_11_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.currState_2_1_LC_2_11_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.dictrl.currState_2_1_LC_2_11_3  (
            .in0(_gnd_net_),
            .in1(N__24673),
            .in2(_gnd_net_),
            .in3(N__20622),
            .lcout(Lab_UT_dictrl_currState_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29406),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_ret_LC_2_11_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_ret_LC_2_11_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.currState_ret_LC_2_11_4 .LUT_INIT=16'b1010111010111111;
    LogicCell40 \Lab_UT.dictrl.currState_ret_LC_2_11_4  (
            .in0(N__24672),
            .in1(N__18061),
            .in2(N__15583),
            .in3(N__14025),
            .lcout(\Lab_UT.dictrl.currState_i_5_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29406),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_fast_0_LC_2_11_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_fast_0_LC_2_11_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.currState_2_fast_0_LC_2_11_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Lab_UT.dictrl.currState_2_fast_0_LC_2_11_5  (
            .in0(_gnd_net_),
            .in1(N__24674),
            .in2(_gnd_net_),
            .in3(N__21109),
            .lcout(\Lab_UT.dictrl.currState_fast_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29406),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_RNITUPT_2_LC_2_11_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_RNITUPT_2_LC_2_11_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_RNITUPT_2_LC_2_11_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Lab_UT.dictrl.currState_2_RNITUPT_2_LC_2_11_6  (
            .in0(N__23344),
            .in1(N__23814),
            .in2(N__25048),
            .in3(N__17887),
            .lcout(\Lab_UT.dictrl.G_30_0_a7_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_3_3_rep1_LC_2_11_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_3_3_rep1_LC_2_11_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.currState_3_3_rep1_LC_2_11_7 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \Lab_UT.dictrl.currState_3_3_rep1_LC_2_11_7  (
            .in0(N__21608),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24675),
            .lcout(\Lab_UT.dictrl.currState_3_rep1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29406),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_0_ret_21_RNIUL8L_0_LC_2_12_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_21_RNIUL8L_0_LC_2_12_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_0_ret_21_RNIUL8L_0_LC_2_12_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_21_RNIUL8L_0_LC_2_12_0  (
            .in0(N__23825),
            .in1(N__18060),
            .in2(_gnd_net_),
            .in3(N__24007),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_11_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_RNIKSEU7_0_0_LC_2_12_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_RNIKSEU7_0_0_LC_2_12_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_RNIKSEU7_0_0_LC_2_12_1 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \Lab_UT.dictrl.currState_2_RNIKSEU7_0_0_LC_2_12_1  (
            .in0(N__21234),
            .in1(N__12313),
            .in2(N__12256),
            .in3(N__27787),
            .lcout(\Lab_UT.dictrl.N_5_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_0_ret_24_LC_2_12_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_24_LC_2_12_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.currState_0_ret_24_LC_2_12_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_24_LC_2_12_2  (
            .in0(N__17567),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15483),
            .lcout(\Lab_UT.dictrl.r_dicLdMtens22_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29399),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_RNIHF8J71_1_LC_2_12_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_RNIHF8J71_1_LC_2_12_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_RNIHF8J71_1_LC_2_12_3 .LUT_INIT=16'b1000110010000000;
    LogicCell40 \Lab_UT.dictrl.currState_2_RNIHF8J71_1_LC_2_12_3  (
            .in0(N__12325),
            .in1(N__21607),
            .in2(N__17892),
            .in3(N__17262),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_RNIDEJTG4_1_LC_2_12_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_RNIDEJTG4_1_LC_2_12_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_RNIDEJTG4_1_LC_2_12_4 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \Lab_UT.dictrl.currState_2_RNIDEJTG4_1_LC_2_12_4  (
            .in0(N__17566),
            .in1(N__15482),
            .in2(N__12319),
            .in3(N__21098),
            .lcout(\Lab_UT.dictrl.N_7_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_3_RNIR9C03_3_LC_2_12_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_3_RNIR9C03_3_LC_2_12_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_3_RNIR9C03_3_LC_2_12_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \Lab_UT.dictrl.currState_3_RNIR9C03_3_LC_2_12_5  (
            .in0(N__18058),
            .in1(N__23824),
            .in2(_gnd_net_),
            .in3(N__27298),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_8_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_ret_5_RNIN6436_0_LC_2_12_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_ret_5_RNIN6436_0_LC_2_12_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_ret_5_RNIN6436_0_LC_2_12_6 .LUT_INIT=16'b1111001011110000;
    LogicCell40 \Lab_UT.dictrl.currState_ret_5_RNIN6436_0_LC_2_12_6  (
            .in0(N__24888),
            .in1(N__18059),
            .in2(N__12316),
            .in3(N__27552),
            .lcout(\Lab_UT.dictrl.N_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_ret_RNI7FNU_LC_2_12_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_ret_RNI7FNU_LC_2_12_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_ret_RNI7FNU_LC_2_12_7 .LUT_INIT=16'b1000100010101010;
    LogicCell40 \Lab_UT.dictrl.currState_ret_RNI7FNU_LC_2_12_7  (
            .in0(N__12307),
            .in1(N__23860),
            .in2(_gnd_net_),
            .in3(N__24889),
            .lcout(\Lab_UT.dictrl.currState_ret_RNI7FNUZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_fast_RNIT3362_0_LC_2_13_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_fast_RNIT3362_0_LC_2_13_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_fast_RNIT3362_0_LC_2_13_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.currState_2_fast_RNIT3362_0_LC_2_13_0  (
            .in0(N__14501),
            .in1(N__17428),
            .in2(N__24901),
            .in3(N__12535),
            .lcout(),
            .ltout(\Lab_UT.dictrl.G_19_0_a7_4_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_fast_RNIOKOT3_0_LC_2_13_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_fast_RNIOKOT3_0_LC_2_13_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_fast_RNIOKOT3_0_LC_2_13_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.currState_2_fast_RNIOKOT3_0_LC_2_13_1  (
            .in0(N__12541),
            .in1(N__18187),
            .in2(N__12301),
            .in3(N__17668),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_0_rep2_RNI0FS1A_LC_2_13_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_0_rep2_RNI0FS1A_LC_2_13_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_0_rep2_RNI0FS1A_LC_2_13_2 .LUT_INIT=16'b1111111111110010;
    LogicCell40 \Lab_UT.dictrl.currState_2_0_rep2_RNI0FS1A_LC_2_13_2  (
            .in0(N__12547),
            .in1(N__24477),
            .in2(N__12298),
            .in3(N__12286),
            .lcout(\Lab_UT.dictrl.G_19_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_ret_5_RNIIF461_LC_2_13_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_ret_5_RNIIF461_LC_2_13_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_ret_5_RNIIF461_LC_2_13_3 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \Lab_UT.dictrl.currState_ret_5_RNIIF461_LC_2_13_3  (
            .in0(N__18057),
            .in1(N__17855),
            .in2(N__24900),
            .in3(N__12295),
            .lcout(\Lab_UT.dictrl.G_19_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_0_rep2_RNI5U4U_LC_2_13_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_0_rep2_RNI5U4U_LC_2_13_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_0_rep2_RNI5U4U_LC_2_13_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.currState_2_0_rep2_RNI5U4U_LC_2_13_5  (
            .in0(N__18056),
            .in1(N__17854),
            .in2(N__20940),
            .in3(N__20369),
            .lcout(\Lab_UT.dictrl.G_19_0_a7_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_6_rep1_RNI4H7E_LC_2_13_6 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_6_rep1_RNI4H7E_LC_2_13_6 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.shifter_6_rep1_RNI4H7E_LC_2_13_6 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \buart.Z_rx.shifter_6_rep1_RNI4H7E_LC_2_13_6  (
            .in0(N__23422),
            .in1(N__22000),
            .in2(N__17910),
            .in3(N__21415),
            .lcout(G_19_0_a7_4_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_4_rep1_RNI7DDT_LC_2_14_6 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_4_rep1_RNI7DDT_LC_2_14_6 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.shifter_4_rep1_RNI7DDT_LC_2_14_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \buart.Z_rx.shifter_4_rep1_RNI7DDT_LC_2_14_6  (
            .in0(_gnd_net_),
            .in1(N__21841),
            .in2(_gnd_net_),
            .in3(N__21444),
            .lcout(G_19_0_a7_4_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.hh_1_LC_2_15_2 .C_ON=1'b0;
    defparam \buart.Z_rx.hh_1_LC_2_15_2 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.hh_1_LC_2_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.hh_1_LC_2_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14292),
            .lcout(\buart.Z_rx.hhZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29383),
            .ce(),
            .sr(N__26087));
    defparam \uu0.l_precount_0_LC_4_1_1 .C_ON=1'b0;
    defparam \uu0.l_precount_0_LC_4_1_1 .SEQ_MODE=4'b1010;
    defparam \uu0.l_precount_0_LC_4_1_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \uu0.l_precount_0_LC_4_1_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12512),
            .lcout(\uu0.l_precountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29470),
            .ce(),
            .sr(N__26093));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_4_2_0 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_4_2_0 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_4_2_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_4_2_0  (
            .in0(_gnd_net_),
            .in1(N__12426),
            .in2(_gnd_net_),
            .in3(N__12373),
            .lcout(\uu0.un99_ci_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_5_LC_4_3_0 .C_ON=1'b0;
    defparam \uu0.l_count_5_LC_4_3_0 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_5_LC_4_3_0 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \uu0.l_count_5_LC_4_3_0  (
            .in0(N__12411),
            .in1(N__12481),
            .in2(_gnd_net_),
            .in3(N__12450),
            .lcout(\uu0.l_countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29455),
            .ce(N__12346),
            .sr(N__26089));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_4_3_2 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_4_3_2 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_4_3_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_4_3_2  (
            .in0(_gnd_net_),
            .in1(N__12480),
            .in2(_gnd_net_),
            .in3(N__12449),
            .lcout(\uu0.un88_ci_3 ),
            .ltout(\uu0.un88_ci_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_6_LC_4_3_3 .C_ON=1'b0;
    defparam \uu0.l_count_6_LC_4_3_3 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_6_LC_4_3_3 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \uu0.l_count_6_LC_4_3_3  (
            .in0(N__12374),
            .in1(N__12412),
            .in2(N__12382),
            .in3(N__13007),
            .lcout(\uu0.l_countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29455),
            .ce(N__12346),
            .sr(N__26089));
    defparam \uu2.mem0.ram512X8_inst_RNO_7_LC_4_3_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_7_LC_4_3_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_7_LC_4_3_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_7_LC_4_3_4  (
            .in0(N__16645),
            .in1(N__16177),
            .in2(_gnd_net_),
            .in3(N__18775),
            .lcout(\uu2.mem0.w_addr_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vram_rd_clk_det_RNI95711_1_LC_4_3_5 .C_ON=1'b0;
    defparam \uu2.vram_rd_clk_det_RNI95711_1_LC_4_3_5 .SEQ_MODE=4'b0000;
    defparam \uu2.vram_rd_clk_det_RNI95711_1_LC_4_3_5 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \uu2.vram_rd_clk_det_RNI95711_1_LC_4_3_5  (
            .in0(N__12625),
            .in1(N__12613),
            .in2(_gnd_net_),
            .in3(N__26144),
            .lcout(\uu2.vram_rd_clk_det_RNI95711Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Mones_subtractor.q20_0_i_LC_4_3_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mones_subtractor.q20_0_i_LC_4_3_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Mones_subtractor.q20_0_i_LC_4_3_6 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \Lab_UT.didp.Mones_subtractor.q20_0_i_LC_4_3_6  (
            .in0(N__26145),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26929),
            .lcout(\Lab_UT.didp.q20_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.uu0.l_count_RNIP43E_13_LC_4_3_7 .C_ON=1'b0;
    defparam \Lab_UT.uu0.l_count_RNIP43E_13_LC_4_3_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.uu0.l_count_RNIP43E_13_LC_4_3_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.uu0.l_count_RNIP43E_13_LC_4_3_7  (
            .in0(_gnd_net_),
            .in1(N__16033),
            .in2(_gnd_net_),
            .in3(N__16009),
            .lcout(\Lab_UT.uu0.un4_l_count_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_12_LC_4_4_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_12_LC_4_4_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_12_LC_4_4_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_12_LC_4_4_0  (
            .in0(N__12666),
            .in1(N__22639),
            .in2(_gnd_net_),
            .in3(N__18798),
            .lcout(\uu2.mem0.w_data_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_13_LC_4_4_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_13_LC_4_4_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_13_LC_4_4_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_13_LC_4_4_1  (
            .in0(N__18799),
            .in1(N__12568),
            .in2(_gnd_net_),
            .in3(N__22618),
            .lcout(\uu2.mem0.w_data_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIOA9K6_8_LC_4_4_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIOA9K6_8_LC_4_4_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIOA9K6_8_LC_4_4_2 .LUT_INIT=16'b1111111100000100;
    LogicCell40 \uu2.w_addr_displaying_RNIOA9K6_8_LC_4_4_2  (
            .in0(N__16399),
            .in1(N__13024),
            .in2(N__16057),
            .in3(N__18864),
            .lcout(\uu2.N_37 ),
            .ltout(\uu2.N_37_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_11_LC_4_4_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_11_LC_4_4_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_11_LC_4_4_3 .LUT_INIT=16'b1101110111011000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_11_LC_4_4_3  (
            .in0(N__18801),
            .in1(N__22834),
            .in2(N__12562),
            .in3(N__12870),
            .lcout(\uu2.mem0.w_data_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_9_LC_4_4_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_9_LC_4_4_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_9_LC_4_4_4 .LUT_INIT=16'b1100110011111010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_9_LC_4_4_4  (
            .in0(N__12667),
            .in1(N__22666),
            .in2(N__12874),
            .in3(N__18802),
            .lcout(\uu2.mem0.w_data_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI7QIF3_8_LC_4_4_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI7QIF3_8_LC_4_4_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI7QIF3_8_LC_4_4_5 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \uu2.w_addr_displaying_RNI7QIF3_8_LC_4_4_5  (
            .in0(N__13023),
            .in1(N__16053),
            .in2(_gnd_net_),
            .in3(N__16398),
            .lcout(),
            .ltout(\uu2.N_51_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIEK5V6_0_LC_4_4_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIEK5V6_0_LC_4_4_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIEK5V6_0_LC_4_4_6 .LUT_INIT=16'b1111000011111100;
    LogicCell40 \uu2.w_addr_displaying_RNIEK5V6_0_LC_4_4_6  (
            .in0(_gnd_net_),
            .in1(N__18865),
            .in2(N__12670),
            .in3(N__19494),
            .lcout(\uu2.N_34 ),
            .ltout(\uu2.N_34_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_8_LC_4_4_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_8_LC_4_4_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_8_LC_4_4_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_8_LC_4_4_7  (
            .in0(N__18800),
            .in1(_gnd_net_),
            .in2(N__12658),
            .in3(N__25682),
            .lcout(\uu2.mem0.w_data_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIASLS1_4_LC_4_5_0 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIASLS1_4_LC_4_5_0 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIASLS1_4_LC_4_5_0 .LUT_INIT=16'b0110010101101010;
    LogicCell40 \uu2.w_addr_displaying_RNIASLS1_4_LC_4_5_0  (
            .in0(N__14919),
            .in1(N__16512),
            .in2(N__14590),
            .in3(N__16275),
            .lcout(),
            .ltout(\uu2.bitmap_pmux_sn_m15_0_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIIO5V6_2_LC_4_5_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIIO5V6_2_LC_4_5_1 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIIO5V6_2_LC_4_5_1 .LUT_INIT=16'b1100101010100000;
    LogicCell40 \uu2.w_addr_displaying_RNIIO5V6_2_LC_4_5_1  (
            .in0(N__12862),
            .in1(N__12646),
            .in2(N__12649),
            .in3(N__14589),
            .lcout(\uu2.bitmap_pmux_sn_i7_mux_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIV2MM2_2_LC_4_5_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIV2MM2_2_LC_4_5_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIV2MM2_2_LC_4_5_2 .LUT_INIT=16'b1000000000010000;
    LogicCell40 \uu2.w_addr_displaying_RNIV2MM2_2_LC_4_5_2  (
            .in0(N__14918),
            .in1(N__19493),
            .in2(N__13525),
            .in3(N__16274),
            .lcout(\uu2.bitmap_pmux_sn_N_65 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI03P31_4_LC_4_5_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI03P31_4_LC_4_5_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI03P31_4_LC_4_5_3 .LUT_INIT=16'b0110011000110011;
    LogicCell40 \uu2.w_addr_displaying_RNI03P31_4_LC_4_5_3  (
            .in0(N__16513),
            .in1(N__14920),
            .in2(_gnd_net_),
            .in3(N__16129),
            .lcout(),
            .ltout(\uu2.bitmap_pmux_sn_m24_0_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIEFIL2_0_LC_4_5_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIEFIL2_0_LC_4_5_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIEFIL2_0_LC_4_5_4 .LUT_INIT=16'b0001100000000110;
    LogicCell40 \uu2.w_addr_displaying_RNIEFIL2_0_LC_4_5_4  (
            .in0(N__14585),
            .in1(N__19492),
            .in2(N__12640),
            .in3(N__16273),
            .lcout(),
            .ltout(\uu2.bitmap_pmux_sn_i5_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI0HFE3_8_LC_4_5_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI0HFE3_8_LC_4_5_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI0HFE3_8_LC_4_5_5 .LUT_INIT=16'b0011000011000000;
    LogicCell40 \uu2.w_addr_displaying_RNI0HFE3_8_LC_4_5_5  (
            .in0(_gnd_net_),
            .in1(N__16787),
            .in2(N__12637),
            .in3(N__16643),
            .lcout(),
            .ltout(\uu2.bitmap_pmux_29_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI649331_8_LC_4_5_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI649331_8_LC_4_5_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI649331_8_LC_4_5_6 .LUT_INIT=16'b1110101001000000;
    LogicCell40 \uu2.w_addr_displaying_RNI649331_8_LC_4_5_6  (
            .in0(N__12883),
            .in1(N__13705),
            .in2(N__12877),
            .in3(N__13501),
            .lcout(\uu2.bitmap_pmux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI12TI1_5_LC_4_5_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI12TI1_5_LC_4_5_7 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI12TI1_5_LC_4_5_7 .LUT_INIT=16'b0010000010100000;
    LogicCell40 \uu2.w_addr_displaying_RNI12TI1_5_LC_4_5_7  (
            .in0(N__16549),
            .in1(N__16786),
            .in2(N__16447),
            .in3(N__16642),
            .lcout(\uu2.bitmap_pmux_sn_N_36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_7_LC_4_6_0 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_7_LC_4_6_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_7_LC_4_6_0 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \buart.Z_tx.shifter_7_LC_4_6_0  (
            .in0(_gnd_net_),
            .in1(N__12830),
            .in2(N__12745),
            .in3(N__12856),
            .lcout(\buart.Z_tx.shifterZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29432),
            .ce(N__12736),
            .sr(N__26082));
    defparam \buart.Z_tx.shifter_8_LC_4_6_1 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_8_LC_4_6_1 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_8_LC_4_6_1 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \buart.Z_tx.shifter_8_LC_4_6_1  (
            .in0(N__12831),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12757),
            .lcout(\buart.Z_tx.shifterZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29432),
            .ce(N__12736),
            .sr(N__26082));
    defparam \uu0.delay_line_RNILLLG7_1_LC_4_6_2 .C_ON=1'b0;
    defparam \uu0.delay_line_RNILLLG7_1_LC_4_6_2 .SEQ_MODE=4'b0000;
    defparam \uu0.delay_line_RNILLLG7_1_LC_4_6_2 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \uu0.delay_line_RNILLLG7_1_LC_4_6_2  (
            .in0(N__12892),
            .in1(N__12915),
            .in2(_gnd_net_),
            .in3(N__13011),
            .lcout(\uu0.un11_l_count_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNIUEOT_58_LC_4_6_3 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIUEOT_58_LC_4_6_3 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIUEOT_58_LC_4_6_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \uu2.bitmap_RNIUEOT_58_LC_4_6_3  (
            .in0(N__16816),
            .in1(N__19084),
            .in2(_gnd_net_),
            .in3(N__16788),
            .lcout(\uu2.N_161 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_6_LC_4_6_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_6_LC_4_6_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_6_LC_4_6_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_6_LC_4_6_4  (
            .in0(N__16789),
            .in1(N__16159),
            .in2(_gnd_net_),
            .in3(N__18786),
            .lcout(\uu2.mem0.w_addr_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_0_LC_4_6_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_0_LC_4_6_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_0_LC_4_6_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_0_LC_4_6_5  (
            .in0(N__16132),
            .in1(N__18973),
            .in2(_gnd_net_),
            .in3(N__18785),
            .lcout(\uu2.mem0.w_addr_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_nesr_RNI4JSO_1_LC_4_6_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_RNI4JSO_1_LC_4_6_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_nesr_RNI4JSO_1_LC_4_6_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.w_addr_displaying_nesr_RNI4JSO_1_LC_4_6_6  (
            .in0(_gnd_net_),
            .in1(N__19487),
            .in2(_gnd_net_),
            .in3(N__16130),
            .lcout(\uu2.N_31_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI25P31_8_LC_4_6_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI25P31_8_LC_4_6_7 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI25P31_8_LC_4_6_7 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \uu2.w_addr_displaying_RNI25P31_8_LC_4_6_7  (
            .in0(N__16131),
            .in1(_gnd_net_),
            .in2(N__19498),
            .in3(N__16644),
            .lcout(\uu2.w_data_displaying_2_i_a2_i_a3_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.sec_clk_LC_4_7_0 .C_ON=1'b0;
    defparam \uu0.sec_clk_LC_4_7_0 .SEQ_MODE=4'b1010;
    defparam \uu0.sec_clk_LC_4_7_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu0.sec_clk_LC_4_7_0  (
            .in0(_gnd_net_),
            .in1(N__26794),
            .in2(_gnd_net_),
            .in3(N__13012),
            .lcout(o_One_Sec_Pulse),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29423),
            .ce(),
            .sr(N__26081));
    defparam \uu2.l_count_1_LC_4_7_1 .C_ON=1'b0;
    defparam \uu2.l_count_1_LC_4_7_1 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_1_LC_4_7_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.l_count_1_LC_4_7_1  (
            .in0(_gnd_net_),
            .in1(N__13078),
            .in2(_gnd_net_),
            .in3(N__13114),
            .lcout(\uu2.l_countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29423),
            .ce(),
            .sr(N__26081));
    defparam \uu2.l_count_0_LC_4_7_2 .C_ON=1'b0;
    defparam \uu2.l_count_0_LC_4_7_2 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_0_LC_4_7_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \uu2.l_count_0_LC_4_7_2  (
            .in0(N__13079),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uu2.l_countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29423),
            .ce(),
            .sr(N__26081));
    defparam \uu2.vram_rd_clk_LC_4_7_3 .C_ON=1'b0;
    defparam \uu2.vram_rd_clk_LC_4_7_3 .SEQ_MODE=4'b1011;
    defparam \uu2.vram_rd_clk_LC_4_7_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.vram_rd_clk_LC_4_7_3  (
            .in0(_gnd_net_),
            .in1(N__13450),
            .in2(_gnd_net_),
            .in3(N__12940),
            .lcout(\uu2.vram_rd_clkZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29423),
            .ce(),
            .sr(N__26081));
    defparam \Lab_UT.uu0.delay_line_1_LC_4_7_4 .C_ON=1'b0;
    defparam \Lab_UT.uu0.delay_line_1_LC_4_7_4 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.uu0.delay_line_1_LC_4_7_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.uu0.delay_line_1_LC_4_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22153),
            .lcout(\Lab_UT.uu0.delay_lineZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29423),
            .ce(),
            .sr(N__26081));
    defparam \uu0.delay_line_1_LC_4_7_7 .C_ON=1'b0;
    defparam \uu0.delay_line_1_LC_4_7_7 .SEQ_MODE=4'b1010;
    defparam \uu0.delay_line_1_LC_4_7_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu0.delay_line_1_LC_4_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12919),
            .lcout(\uu0.delay_lineZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29423),
            .ce(),
            .sr(N__26081));
    defparam \Lab_UT.dictrl.currState_ret_2_LC_4_8_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_ret_2_LC_4_8_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.currState_ret_2_LC_4_8_1 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \Lab_UT.dictrl.currState_ret_2_LC_4_8_1  (
            .in0(N__24626),
            .in1(N__20814),
            .in2(_gnd_net_),
            .in3(N__21624),
            .lcout(\Lab_UT.dictrl.r_dicLdMtens23_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29414),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_0_LC_4_8_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_0_LC_4_8_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.currState_2_0_LC_4_8_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Lab_UT.dictrl.currState_2_0_LC_4_8_2  (
            .in0(_gnd_net_),
            .in1(N__24627),
            .in2(_gnd_net_),
            .in3(N__21108),
            .lcout(\Lab_UT.dictrl.currStateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29414),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.sec_clkD_RNISDHD_LC_4_8_3 .C_ON=1'b0;
    defparam \uu0.sec_clkD_RNISDHD_LC_4_8_3 .SEQ_MODE=4'b0000;
    defparam \uu0.sec_clkD_RNISDHD_LC_4_8_3 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \uu0.sec_clkD_RNISDHD_LC_4_8_3  (
            .in0(N__26784),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26748),
            .lcout(oneSecStrb),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.sec_clkD_LC_4_8_4 .C_ON=1'b0;
    defparam \uu0.sec_clkD_LC_4_8_4 .SEQ_MODE=4'b1000;
    defparam \uu0.sec_clkD_LC_4_8_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu0.sec_clkD_LC_4_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26785),
            .lcout(uu0_sec_clkD),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29414),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_count.counter_gen_label_2__un284_ci_LC_4_8_5 .C_ON=1'b0;
    defparam \uu2.vbuf_count.counter_gen_label_2__un284_ci_LC_4_8_5 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_count.counter_gen_label_2__un284_ci_LC_4_8_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.vbuf_count.counter_gen_label_2__un284_ci_LC_4_8_5  (
            .in0(_gnd_net_),
            .in1(N__13113),
            .in2(_gnd_net_),
            .in3(N__13077),
            .lcout(\uu2.un284_ci ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_ness_RNO_0_6_LC_4_8_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_ness_RNO_0_6_LC_4_8_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_ness_RNO_0_6_LC_4_8_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \uu2.w_addr_displaying_ness_RNO_0_6_LC_4_8_6  (
            .in0(_gnd_net_),
            .in1(N__16465),
            .in2(_gnd_net_),
            .in3(N__16375),
            .lcout(\uu2.N_48 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.rst_LC_4_9_0 .C_ON=1'b0;
    defparam \resetGen.rst_LC_4_9_0 .SEQ_MODE=4'b1000;
    defparam \resetGen.rst_LC_4_9_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \resetGen.rst_LC_4_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19191),
            .lcout(rst),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29407),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_ret_RNI5RB74_LC_4_9_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_ret_RNI5RB74_LC_4_9_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_ret_RNI5RB74_LC_4_9_1 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \Lab_UT.dictrl.currState_ret_RNI5RB74_LC_4_9_1  (
            .in0(N__27295),
            .in1(N__13896),
            .in2(_gnd_net_),
            .in3(N__27792),
            .lcout(\Lab_UT.dictrl.dicLdAMtens_rst ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__m8_LC_4_9_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__m8_LC_4_9_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__m8_LC_4_9_2 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__m8_LC_4_9_2  (
            .in0(N__20392),
            .in1(N__14179),
            .in2(_gnd_net_),
            .in3(N__14161),
            .lcout(\Lab_UT.dictrl.N_9 ),
            .ltout(\Lab_UT.dictrl.N_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_RNINHPTJ_1_LC_4_9_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_RNINHPTJ_1_LC_4_9_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_RNINHPTJ_1_LC_4_9_3 .LUT_INIT=16'b1000000010100010;
    LogicCell40 \Lab_UT.dictrl.currState_2_RNINHPTJ_1_LC_4_9_3  (
            .in0(N__13948),
            .in1(N__17916),
            .in2(N__13030),
            .in3(N__20284),
            .lcout(\Lab_UT.dictrl.N_19_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_RNIR9C03_2_LC_4_9_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_RNIR9C03_2_LC_4_9_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_RNIR9C03_2_LC_4_9_4 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \Lab_UT.dictrl.currState_2_RNIR9C03_2_LC_4_9_4  (
            .in0(N__25008),
            .in1(N__23430),
            .in2(N__23833),
            .in3(N__27294),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_21_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_ret_5_RNIN6436_LC_4_9_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_ret_5_RNIN6436_LC_4_9_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_ret_5_RNIN6436_LC_4_9_5 .LUT_INIT=16'b1111001011110000;
    LogicCell40 \Lab_UT.dictrl.currState_ret_5_RNIN6436_LC_4_9_5  (
            .in0(N__24864),
            .in1(N__18014),
            .in2(N__13027),
            .in3(N__27551),
            .lcout(\Lab_UT.dictrl.N_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_0_0_LC_4_9_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_0_0_LC_4_9_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_0_0_LC_4_9_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__g0_0_0_LC_4_9_6  (
            .in0(_gnd_net_),
            .in1(N__14101),
            .in2(_gnd_net_),
            .in3(N__27293),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_1_LC_4_9_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_1_LC_4_9_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_1_LC_4_9_7 .LUT_INIT=16'b1011100010001000;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__g0_1_LC_4_9_7  (
            .in0(N__23972),
            .in1(N__23827),
            .in2(N__13138),
            .in3(N__27791),
            .lcout(\Lab_UT.dictrl.N_23_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__m21_mb_LC_4_10_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__m21_mb_LC_4_10_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__m21_mb_LC_4_10_0 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__m21_mb_LC_4_10_0  (
            .in0(N__13144),
            .in1(N__23818),
            .in2(N__25039),
            .in3(N__14455),
            .lcout(\Lab_UT.dictrl.i8_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_0_ret_21_LC_4_10_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_21_LC_4_10_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.currState_0_ret_21_LC_4_10_1 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_21_LC_4_10_1  (
            .in0(N__13192),
            .in1(N__13183),
            .in2(N__13126),
            .in3(N__13168),
            .lcout(\Lab_UT.dictrl.currState_i_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29400),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_0_ret_1_RNINTRN4_LC_4_10_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_1_RNINTRN4_LC_4_10_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_0_ret_1_RNINTRN4_LC_4_10_2 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_1_RNINTRN4_LC_4_10_2  (
            .in0(N__27747),
            .in1(N__23898),
            .in2(_gnd_net_),
            .in3(N__27277),
            .lcout(\Lab_UT.dictrl.dicLdAStens_rst ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_RNIA8EV3_0_1_LC_4_10_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_RNIA8EV3_0_1_LC_4_10_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_RNIA8EV3_0_1_LC_4_10_3 .LUT_INIT=16'b1110010011110101;
    LogicCell40 \Lab_UT.dictrl.nextState_RNIA8EV3_0_1_LC_4_10_3  (
            .in0(N__23381),
            .in1(N__13252),
            .in2(N__13237),
            .in3(N__27745),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_1611_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_RNIFHD18_1_LC_4_10_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_RNIFHD18_1_LC_4_10_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_RNIFHD18_1_LC_4_10_4 .LUT_INIT=16'b0011000011111100;
    LogicCell40 \Lab_UT.dictrl.nextState_RNIFHD18_1_LC_4_10_4  (
            .in0(_gnd_net_),
            .in1(N__18006),
            .in2(N__13135),
            .in3(N__13132),
            .lcout(\Lab_UT.dictrl.N_1605_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_3_RNI3HN91_3_LC_4_10_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_3_RNI3HN91_3_LC_4_10_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_3_RNI3HN91_3_LC_4_10_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \Lab_UT.dictrl.currState_3_RNI3HN91_3_LC_4_10_5  (
            .in0(N__14209),
            .in1(N__23817),
            .in2(_gnd_net_),
            .in3(N__18115),
            .lcout(\Lab_UT.dictrl.G_28_0_a5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_RNI0LLB7_0_LC_4_10_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_RNI0LLB7_0_LC_4_10_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_RNI0LLB7_0_LC_4_10_6 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \Lab_UT.dictrl.currState_2_RNI0LLB7_0_LC_4_10_6  (
            .in0(N__27746),
            .in1(N__15349),
            .in2(N__21244),
            .in3(N__27276),
            .lcout(\Lab_UT.dictrl.N_8_3 ),
            .ltout(\Lab_UT.dictrl.N_8_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_RNIQ7IPD1_0_LC_4_10_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_RNIQ7IPD1_0_LC_4_10_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_RNIQ7IPD1_0_LC_4_10_7 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \Lab_UT.dictrl.currState_2_RNIQ7IPD1_0_LC_4_10_7  (
            .in0(N__13191),
            .in1(N__13182),
            .in2(N__13174),
            .in3(N__13167),
            .lcout(\Lab_UT.dictrl.N_6ctr ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_0_rep2_RNIBGCI9_LC_4_11_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_0_rep2_RNIBGCI9_LC_4_11_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_0_rep2_RNIBGCI9_LC_4_11_0 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \Lab_UT.dictrl.currState_2_0_rep2_RNIBGCI9_LC_4_11_0  (
            .in0(N__13153),
            .in1(N__14107),
            .in2(N__13279),
            .in3(N__13159),
            .lcout(),
            .ltout(\Lab_UT.dictrl.currState_2_0_rep2_RNIBGCIZ0Z9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_RNI0GB6H_0_LC_4_11_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_RNI0GB6H_0_LC_4_11_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_RNI0GB6H_0_LC_4_11_1 .LUT_INIT=16'b1000000011000100;
    LogicCell40 \Lab_UT.dictrl.nextState_RNI0GB6H_0_LC_4_11_1  (
            .in0(N__18111),
            .in1(N__14205),
            .in2(N__13171),
            .in3(N__13981),
            .lcout(\Lab_UT.dictrl.G_28_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_0_rep2_RNIKH8P2_LC_4_11_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_0_rep2_RNIKH8P2_LC_4_11_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_0_rep2_RNIKH8P2_LC_4_11_2 .LUT_INIT=16'b0001000100110011;
    LogicCell40 \Lab_UT.dictrl.currState_2_0_rep2_RNIKH8P2_LC_4_11_2  (
            .in0(N__20936),
            .in1(N__29073),
            .in2(_gnd_net_),
            .in3(N__27248),
            .lcout(\Lab_UT.dictrl.currState_2_0_rep2_RNIKH8PZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_RNI0KKK6_0_LC_4_11_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_RNI0KKK6_0_LC_4_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_RNI0KKK6_0_LC_4_11_3 .LUT_INIT=16'b1111101001110010;
    LogicCell40 \Lab_UT.dictrl.nextState_RNI0KKK6_0_LC_4_11_3  (
            .in0(N__18041),
            .in1(N__24813),
            .in2(N__14008),
            .in3(N__13243),
            .lcout(\Lab_UT.dictrl.N_1609_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_RNIS6CF1_5_LC_4_11_4 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_RNIS6CF1_5_LC_4_11_4 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.shifter_RNIS6CF1_5_LC_4_11_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \buart.Z_rx.shifter_RNIS6CF1_5_LC_4_11_4  (
            .in0(N__28981),
            .in1(N__24448),
            .in2(_gnd_net_),
            .in3(N__27731),
            .lcout(shifter_RNIS6CF1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_4_LC_4_11_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_4_LC_4_11_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_4_LC_4_11_5 .LUT_INIT=16'b0010110011101100;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__g0_4_LC_4_11_5  (
            .in0(N__27247),
            .in1(N__20937),
            .in2(N__27788),
            .in3(N__27517),
            .lcout(\Lab_UT.dictrl.N_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__m21_rn_1_0_LC_4_11_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__m21_rn_1_0_LC_4_11_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__m21_rn_1_0_LC_4_11_6 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__m21_rn_1_0_LC_4_11_6  (
            .in0(N__20935),
            .in1(N__27730),
            .in2(_gnd_net_),
            .in3(N__27249),
            .lcout(),
            .ltout(\Lab_UT.dictrl.m21_rn_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__m21_rn_LC_4_11_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__m21_rn_LC_4_11_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__m21_rn_LC_4_11_7 .LUT_INIT=16'b0111001011111010;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__m21_rn_LC_4_11_7  (
            .in0(N__25012),
            .in1(N__24814),
            .in2(N__13147),
            .in3(N__15320),
            .lcout(\Lab_UT.dictrl.m21_rn_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_ret_5_LC_4_12_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_ret_5_LC_4_12_0 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.currState_ret_5_LC_4_12_0 .LUT_INIT=16'b0001101110111011;
    LogicCell40 \Lab_UT.dictrl.currState_ret_5_LC_4_12_0  (
            .in0(N__18046),
            .in1(N__13957),
            .in2(N__13974),
            .in3(N__17915),
            .lcout(\Lab_UT.dictrl.currState_i_5_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29389),
            .ce(),
            .sr(N__26064));
    defparam \Lab_UT.dictrl.currState_2_0_rep1_RNI3BNS2_LC_4_12_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_0_rep1_RNI3BNS2_LC_4_12_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_0_rep1_RNI3BNS2_LC_4_12_1 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \Lab_UT.dictrl.currState_2_0_rep1_RNI3BNS2_LC_4_12_1  (
            .in0(N__27483),
            .in1(N__24802),
            .in2(_gnd_net_),
            .in3(N__14088),
            .lcout(\Lab_UT.dictrl.g1_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_17_LC_4_12_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_17_LC_4_12_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_17_LC_4_12_2 .LUT_INIT=16'b0101110011111100;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__g0_17_LC_4_12_2  (
            .in0(N__27645),
            .in1(N__14347),
            .in2(N__14096),
            .in3(N__27212),
            .lcout(\Lab_UT.dictrl.N_13_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_18_LC_4_12_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_18_LC_4_12_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_18_LC_4_12_3 .LUT_INIT=16'b0010111011001100;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__g0_18_LC_4_12_3  (
            .in0(N__27210),
            .in1(N__14087),
            .in2(N__27510),
            .in3(N__27646),
            .lcout(\Lab_UT.dictrl.N_7_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__m4_LC_4_12_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__m4_LC_4_12_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__m4_LC_4_12_4 .LUT_INIT=16'b0101100011111000;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__m4_LC_4_12_4  (
            .in0(N__27643),
            .in1(N__27475),
            .in2(N__14095),
            .in3(N__27209),
            .lcout(\Lab_UT.dictrl.N_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__m6_LC_4_12_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__m6_LC_4_12_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__m6_LC_4_12_5 .LUT_INIT=16'b0010111011001100;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__m6_LC_4_12_5  (
            .in0(N__27211),
            .in1(N__14083),
            .in2(N__27511),
            .in3(N__27644),
            .lcout(\Lab_UT.dictrl.N_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__m19_LC_4_12_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__m19_LC_4_12_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__m19_LC_4_12_6 .LUT_INIT=16'b1000000010000000;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__m19_LC_4_12_6  (
            .in0(N__27647),
            .in1(N__27482),
            .in2(N__14097),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.dictrl.N_20 ),
            .ltout(\Lab_UT.dictrl.N_20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_RNIA8EV3_1_LC_4_12_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_RNIA8EV3_1_LC_4_12_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_RNIA8EV3_1_LC_4_12_7 .LUT_INIT=16'b1010101000111111;
    LogicCell40 \Lab_UT.dictrl.nextState_RNIA8EV3_1_LC_4_12_7  (
            .in0(N__13233),
            .in1(N__24803),
            .in2(N__13195),
            .in3(N__23431),
            .lcout(\Lab_UT.dictrl.nextState_RNIA8EV3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.decoder.de_littleA_2_0_LC_4_13_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.decoder.de_littleA_2_0_LC_4_13_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.decoder.de_littleA_2_0_LC_4_13_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Lab_UT.dictrl.decoder.de_littleA_2_0_LC_4_13_0  (
            .in0(N__21389),
            .in1(N__21441),
            .in2(N__21767),
            .in3(N__21683),
            .lcout(\Lab_UT.dictrl.decoder.de_littleA_2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.decoder.de_num_0_LC_4_13_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.decoder.de_num_0_LC_4_13_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.decoder.de_num_0_LC_4_13_1 .LUT_INIT=16'b0010001000101010;
    LogicCell40 \Lab_UT.dictrl.decoder.de_num_0_LC_4_13_1  (
            .in0(N__14223),
            .in1(N__21749),
            .in2(N__21698),
            .in3(N__21392),
            .lcout(\Lab_UT.dictrl.de_num_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.decoder.de_num0to5_1_LC_4_13_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.decoder.de_num0to5_1_LC_4_13_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.decoder.de_num0to5_1_LC_4_13_2 .LUT_INIT=16'b0000011100000000;
    LogicCell40 \Lab_UT.dictrl.decoder.de_num0to5_1_LC_4_13_2  (
            .in0(N__21391),
            .in1(N__21685),
            .in2(N__21766),
            .in3(N__14222),
            .lcout(\Lab_UT.dictrl.de_num0to5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.decoder.g0_1_LC_4_13_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.decoder.g0_1_LC_4_13_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.decoder.g0_1_LC_4_13_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Lab_UT.dictrl.decoder.g0_1_LC_4_13_3  (
            .in0(_gnd_net_),
            .in1(N__21390),
            .in2(_gnd_net_),
            .in3(N__21352),
            .lcout(\Lab_UT.dictrl.decoder.g0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.decoder.g0_5_LC_4_13_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.decoder.g0_5_LC_4_13_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.decoder.g0_5_LC_4_13_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.decoder.g0_5_LC_4_13_4  (
            .in0(N__21756),
            .in1(N__21684),
            .in2(N__21999),
            .in3(N__21936),
            .lcout(),
            .ltout(\Lab_UT.dictrl.decoder.g0Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.decoder.g0_6_LC_4_13_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.decoder.g0_6_LC_4_13_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.decoder.g0_6_LC_4_13_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Lab_UT.dictrl.decoder.g0_6_LC_4_13_5  (
            .in0(N__25372),
            .in1(N__25272),
            .in2(N__13264),
            .in3(N__13261),
            .lcout(\Lab_UT.dictrl.g0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_21_LC_4_13_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_21_LC_4_13_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_21_LC_4_13_6 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__g0_21_LC_4_13_6  (
            .in0(N__21222),
            .in1(N__27773),
            .in2(N__18400),
            .in3(N__27246),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_36_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_20_LC_4_13_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_20_LC_4_13_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_20_LC_4_13_7 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__g0_20_LC_4_13_7  (
            .in0(N__14239),
            .in1(N__15304),
            .in2(N__13255),
            .in3(N__23815),
            .lcout(\Lab_UT.dictrl.N_38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_4_rep1_LC_4_14_0 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_4_rep1_LC_4_14_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_4_rep1_LC_4_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_4_rep1_LC_4_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24415),
            .lcout(bu_rx_data_4_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29380),
            .ce(N__25428),
            .sr(N__26090));
    defparam \buart.Z_rx.shifter_1_rep1_LC_4_14_1 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_1_rep1_LC_4_14_1 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_1_rep1_LC_4_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_1_rep1_LC_4_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28596),
            .lcout(bu_rx_data_1_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29380),
            .ce(N__25428),
            .sr(N__26090));
    defparam \buart.Z_rx.shifter_3_rep1_LC_4_14_2 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_3_rep1_LC_4_14_2 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_3_rep1_LC_4_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_3_rep1_LC_4_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25279),
            .lcout(bu_rx_data_3_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29380),
            .ce(N__25428),
            .sr(N__26090));
    defparam \buart.Z_rx.shifter_fast_7_LC_4_14_3 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_7_LC_4_14_3 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_fast_7_LC_4_14_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_fast_7_LC_4_14_3  (
            .in0(N__21877),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_fast_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29380),
            .ce(N__25428),
            .sr(N__26090));
    defparam \buart.Z_rx.shifter_4_LC_4_14_5 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_4_LC_4_14_5 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_4_LC_4_14_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_4_LC_4_14_5  (
            .in0(N__24416),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29380),
            .ce(N__25428),
            .sr(N__26090));
    defparam \buart.Z_rx.shifter_2_rep1_LC_4_14_6 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_2_rep1_LC_4_14_6 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_2_rep1_LC_4_14_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_2_rep1_LC_4_14_6  (
            .in0(N__28982),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_2_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29380),
            .ce(N__25428),
            .sr(N__26090));
    defparam \Lab_UT.dictrl.nextState_1_3_0__m7_LC_4_15_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__m7_LC_4_15_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__m7_LC_4_15_0 .LUT_INIT=16'b1111010011111100;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__m7_LC_4_15_0  (
            .in0(N__27716),
            .in1(N__24004),
            .in2(N__14437),
            .in3(N__14224),
            .lcout(\Lab_UT.dictrl.N_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_3_3_rep1_RNIM4AP_LC_4_15_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_3_3_rep1_RNIM4AP_LC_4_15_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_3_3_rep1_RNIM4AP_LC_4_15_2 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \Lab_UT.dictrl.currState_3_3_rep1_RNIM4AP_LC_4_15_2  (
            .in0(N__25344),
            .in1(N__28613),
            .in2(_gnd_net_),
            .in3(N__20370),
            .lcout(),
            .ltout(G_28_0_a5_0_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_RNI1D8L1_4_LC_4_15_3 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_RNI1D8L1_4_LC_4_15_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.shifter_RNI1D8L1_4_LC_4_15_3 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \buart.Z_rx.shifter_RNI1D8L1_4_LC_4_15_3  (
            .in0(N__28817),
            .in1(N__24266),
            .in2(N__13282),
            .in3(N__25273),
            .lcout(shifter_RNI1D8L1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_6_LC_4_15_4 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_6_LC_4_15_4 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_6_LC_4_15_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_6_LC_4_15_4  (
            .in0(N__25345),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29375),
            .ce(N__25425),
            .sr(N__26092));
    defparam \buart.Z_rx.shifter_fast_6_LC_4_15_6 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_6_LC_4_15_6 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_fast_6_LC_4_15_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_fast_6_LC_4_15_6  (
            .in0(N__25346),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_fast_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29375),
            .ce(N__25425),
            .sr(N__26092));
    defparam \buart.Z_rx.shifter_7_LC_4_15_7 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_7_LC_4_15_7 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_7_LC_4_15_7 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \buart.Z_rx.shifter_7_LC_4_15_7  (
            .in0(_gnd_net_),
            .in1(N__21871),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29375),
            .ce(N__25425),
            .sr(N__26092));
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_4_16_0 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_4_16_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_4_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_4_16_0  (
            .in0(_gnd_net_),
            .in1(N__14415),
            .in2(N__13297),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_16_0_),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_4_16_1 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_4_16_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_4_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_4_16_1  (
            .in0(_gnd_net_),
            .in1(N__13308),
            .in2(_gnd_net_),
            .in3(N__13267),
            .lcout(\buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.Z_baudgen.un5_counter_cry_1 ),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_3_LC_4_16_2 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.counter_3_LC_4_16_2 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_3_LC_4_16_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_3_LC_4_16_2  (
            .in0(N__15926),
            .in1(N__14428),
            .in2(_gnd_net_),
            .in3(N__13339),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_3 ),
            .ltout(),
            .carryin(\buart.Z_rx.Z_baudgen.un5_counter_cry_2 ),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_3 ),
            .clk(N__29373),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_4_16_3 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_4_16_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_4_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_4_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14380),
            .in3(N__13336),
            .lcout(\buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.Z_baudgen.un5_counter_cry_3 ),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_5_LC_4_16_4 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_5_LC_4_16_4 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_5_LC_4_16_4 .LUT_INIT=16'b0000000100000100;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_5_LC_4_16_4  (
            .in0(N__15925),
            .in1(N__13329),
            .in2(N__15625),
            .in3(N__13333),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29373),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_RNI4IE3_5_LC_4_16_5 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI4IE3_5_LC_4_16_5 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI4IE3_5_LC_4_16_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_RNI4IE3_5_LC_4_16_5  (
            .in0(N__14375),
            .in1(N__13307),
            .in2(N__13330),
            .in3(N__13292),
            .lcout(\buart.Z_rx.Z_baudgen.ser_clk_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_2_LC_4_16_6 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_2_LC_4_16_6 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_2_LC_4_16_6 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_2_LC_4_16_6  (
            .in0(N__13309),
            .in1(N__15924),
            .in2(N__13318),
            .in3(N__15624),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29373),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_1_LC_4_16_7 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_1_LC_4_16_7 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_1_LC_4_16_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_1_LC_4_16_7  (
            .in0(N__15923),
            .in1(N__14416),
            .in2(_gnd_net_),
            .in3(N__13296),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29373),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_addr_2_LC_5_3_0 .C_ON=1'b0;
    defparam \uu2.r_addr_2_LC_5_3_0 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_2_LC_5_3_0 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.r_addr_2_LC_5_3_0  (
            .in0(N__13626),
            .in1(N__13589),
            .in2(N__13662),
            .in3(N__25133),
            .lcout(\uu2.r_addrZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29447),
            .ce(),
            .sr(N__26068));
    defparam \uu2.r_addr_1_LC_5_3_1 .C_ON=1'b0;
    defparam \uu2.r_addr_1_LC_5_3_1 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_1_LC_5_3_1 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \uu2.r_addr_1_LC_5_3_1  (
            .in0(N__25132),
            .in1(_gnd_net_),
            .in2(N__13593),
            .in3(N__13625),
            .lcout(\uu2.r_addrZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29447),
            .ce(),
            .sr(N__26068));
    defparam \uu2.trig_rd_det_RNINBDQ_1_LC_5_3_2 .C_ON=1'b0;
    defparam \uu2.trig_rd_det_RNINBDQ_1_LC_5_3_2 .SEQ_MODE=4'b0000;
    defparam \uu2.trig_rd_det_RNINBDQ_1_LC_5_3_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \uu2.trig_rd_det_RNINBDQ_1_LC_5_3_2  (
            .in0(_gnd_net_),
            .in1(N__25131),
            .in2(_gnd_net_),
            .in3(N__26150),
            .lcout(\uu2.trig_rd_is_det_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.trig_rd_det_RNIJIIO_1_LC_5_3_3 .C_ON=1'b0;
    defparam \uu2.trig_rd_det_RNIJIIO_1_LC_5_3_3 .SEQ_MODE=4'b0000;
    defparam \uu2.trig_rd_det_RNIJIIO_1_LC_5_3_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uu2.trig_rd_det_RNIJIIO_1_LC_5_3_3  (
            .in0(_gnd_net_),
            .in1(N__13474),
            .in2(_gnd_net_),
            .in3(N__13407),
            .lcout(\uu2.trig_rd_is_det ),
            .ltout(\uu2.trig_rd_is_det_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_addr_0_LC_5_3_4 .C_ON=1'b0;
    defparam \uu2.r_addr_0_LC_5_3_4 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_0_LC_5_3_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \uu2.r_addr_0_LC_5_3_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13477),
            .in3(N__13585),
            .lcout(\uu2.r_addrZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29447),
            .ce(),
            .sr(N__26068));
    defparam \uu2.trig_rd_det_1_LC_5_3_5 .C_ON=1'b0;
    defparam \uu2.trig_rd_det_1_LC_5_3_5 .SEQ_MODE=4'b1000;
    defparam \uu2.trig_rd_det_1_LC_5_3_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.trig_rd_det_1_LC_5_3_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13408),
            .lcout(\uu2.trig_rd_detZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29447),
            .ce(),
            .sr(N__26068));
    defparam \uu2.trig_rd_det_0_LC_5_3_6 .C_ON=1'b0;
    defparam \uu2.trig_rd_det_0_LC_5_3_6 .SEQ_MODE=4'b1000;
    defparam \uu2.trig_rd_det_0_LC_5_3_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uu2.trig_rd_det_0_LC_5_3_6  (
            .in0(_gnd_net_),
            .in1(N__13467),
            .in2(_gnd_net_),
            .in3(N__13426),
            .lcout(\uu2.trig_rd_detZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29447),
            .ce(),
            .sr(N__26068));
    defparam \uu2.vbuf_raddr.counter_gen_label_8__un448_ci_0_LC_5_4_0 .C_ON=1'b0;
    defparam \uu2.vbuf_raddr.counter_gen_label_8__un448_ci_0_LC_5_4_0 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_raddr.counter_gen_label_8__un448_ci_0_LC_5_4_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.vbuf_raddr.counter_gen_label_8__un448_ci_0_LC_5_4_0  (
            .in0(_gnd_net_),
            .in1(N__13355),
            .in2(_gnd_net_),
            .in3(N__13684),
            .lcout(\uu2.vbuf_raddr.un448_ci_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_raddr.counter_gen_label_6__un426_ci_3_LC_5_4_1 .C_ON=1'b0;
    defparam \uu2.vbuf_raddr.counter_gen_label_6__un426_ci_3_LC_5_4_1 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_raddr.counter_gen_label_6__un426_ci_3_LC_5_4_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uu2.vbuf_raddr.counter_gen_label_6__un426_ci_3_LC_5_4_1  (
            .in0(N__22793),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25109),
            .lcout(\uu2.vbuf_raddr.un426_ci_3 ),
            .ltout(\uu2.vbuf_raddr.un426_ci_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_addr_esr_8_LC_5_4_2 .C_ON=1'b0;
    defparam \uu2.r_addr_esr_8_LC_5_4_2 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_esr_8_LC_5_4_2 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \uu2.r_addr_esr_8_LC_5_4_2  (
            .in0(N__13383),
            .in1(N__13399),
            .in2(N__13393),
            .in3(N__25160),
            .lcout(\uu2.r_addrZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29439),
            .ce(N__13534),
            .sr(N__26066));
    defparam \uu2.r_addr_esr_7_LC_5_4_3 .C_ON=1'b0;
    defparam \uu2.r_addr_esr_7_LC_5_4_3 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_esr_7_LC_5_4_3 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu2.r_addr_esr_7_LC_5_4_3  (
            .in0(N__25161),
            .in1(N__13356),
            .in2(N__13692),
            .in3(N__13369),
            .lcout(\uu2.r_addrZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29439),
            .ce(N__13534),
            .sr(N__26066));
    defparam \uu2.vbuf_raddr.counter_gen_label_4__un404_ci_LC_5_4_4 .C_ON=1'b0;
    defparam \uu2.vbuf_raddr.counter_gen_label_4__un404_ci_LC_5_4_4 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_raddr.counter_gen_label_4__un404_ci_LC_5_4_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.vbuf_raddr.counter_gen_label_4__un404_ci_LC_5_4_4  (
            .in0(N__13654),
            .in1(N__13623),
            .in2(N__13556),
            .in3(N__13583),
            .lcout(\uu2.un404_ci_0 ),
            .ltout(\uu2.un404_ci_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_addr_esr_6_LC_5_4_5 .C_ON=1'b0;
    defparam \uu2.r_addr_esr_6_LC_5_4_5 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_esr_6_LC_5_4_5 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \uu2.r_addr_esr_6_LC_5_4_5  (
            .in0(N__13688),
            .in1(N__22807),
            .in2(N__13699),
            .in3(N__25110),
            .lcout(\uu2.r_addrZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29439),
            .ce(N__13534),
            .sr(N__26066));
    defparam \uu2.r_addr_esr_3_LC_5_4_6 .C_ON=1'b0;
    defparam \uu2.r_addr_esr_3_LC_5_4_6 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_esr_3_LC_5_4_6 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.r_addr_esr_3_LC_5_4_6  (
            .in0(N__13655),
            .in1(N__13624),
            .in2(N__13557),
            .in3(N__13584),
            .lcout(\uu2.r_addrZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29439),
            .ce(N__13534),
            .sr(N__26066));
    defparam \uu2.w_addr_displaying_RNI12TI1_0_5_LC_5_4_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI12TI1_0_5_LC_5_4_7 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI12TI1_0_5_LC_5_4_7 .LUT_INIT=16'b0000001101001000;
    LogicCell40 \uu2.w_addr_displaying_RNI12TI1_0_5_LC_5_4_7  (
            .in0(N__16545),
            .in1(N__16768),
            .in2(N__16442),
            .in3(N__16627),
            .lcout(\uu2.bitmap_pmux_sn_N_42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNIHNN91_40_LC_5_5_0 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIHNN91_40_LC_5_5_0 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIHNN91_40_LC_5_5_0 .LUT_INIT=16'b0000110001110111;
    LogicCell40 \uu2.bitmap_RNIHNN91_40_LC_5_5_0  (
            .in0(N__13762),
            .in1(N__16257),
            .in2(N__13756),
            .in3(N__16640),
            .lcout(),
            .ltout(\uu2.bitmap_pmux_26_bm_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNI1PH82_34_LC_5_5_1 .C_ON=1'b0;
    defparam \uu2.bitmap_RNI1PH82_34_LC_5_5_1 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNI1PH82_34_LC_5_5_1 .LUT_INIT=16'b0101111000001110;
    LogicCell40 \uu2.bitmap_RNI1PH82_34_LC_5_5_1  (
            .in0(N__16258),
            .in1(N__13483),
            .in2(N__13516),
            .in3(N__14950),
            .lcout(\uu2.bitmap_RNI1PH82Z0Z_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI2NHS5_8_LC_5_5_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI2NHS5_8_LC_5_5_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI2NHS5_8_LC_5_5_2 .LUT_INIT=16'b0010000011111101;
    LogicCell40 \uu2.w_addr_displaying_RNI2NHS5_8_LC_5_5_2  (
            .in0(N__16259),
            .in1(N__16641),
            .in2(N__13513),
            .in3(N__14632),
            .lcout(),
            .ltout(\uu2.N_400_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIB4NVD_4_LC_5_5_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIB4NVD_4_LC_5_5_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIB4NVD_4_LC_5_5_3 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \uu2.w_addr_displaying_RNIB4NVD_4_LC_5_5_3  (
            .in0(_gnd_net_),
            .in1(N__14626),
            .in2(N__13504),
            .in3(N__13489),
            .lcout(\uu2.N_409 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNIPUBH6_34_LC_5_5_4 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIPUBH6_34_LC_5_5_4 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIPUBH6_34_LC_5_5_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \uu2.bitmap_RNIPUBH6_34_LC_5_5_4  (
            .in0(N__14929),
            .in1(N__13495),
            .in2(_gnd_net_),
            .in3(N__14608),
            .lcout(\uu2.N_404 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_290_LC_5_5_5 .C_ON=1'b0;
    defparam \uu2.bitmap_290_LC_5_5_5 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_290_LC_5_5_5 .LUT_INIT=16'b1011101010101010;
    LogicCell40 \uu2.bitmap_290_LC_5_5_5  (
            .in0(N__19888),
            .in1(N__17056),
            .in2(N__15064),
            .in3(N__16870),
            .lcout(\uu2.bitmapZ0Z_290 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_290C_net ),
            .ce(),
            .sr(N__26041));
    defparam \uu2.bitmap_40_LC_5_5_6 .C_ON=1'b0;
    defparam \uu2.bitmap_40_LC_5_5_6 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_40_LC_5_5_6 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \uu2.bitmap_40_LC_5_5_6  (
            .in0(N__15118),
            .in1(N__19889),
            .in2(_gnd_net_),
            .in3(N__14863),
            .lcout(\uu2.bitmapZ0Z_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_290C_net ),
            .ce(),
            .sr(N__26041));
    defparam \uu2.bitmap_296_LC_5_5_7 .C_ON=1'b0;
    defparam \uu2.bitmap_296_LC_5_5_7 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_296_LC_5_5_7 .LUT_INIT=16'b1111101011110000;
    LogicCell40 \uu2.bitmap_296_LC_5_5_7  (
            .in0(N__14854),
            .in1(_gnd_net_),
            .in2(N__19897),
            .in3(N__15117),
            .lcout(\uu2.bitmapZ0Z_296 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_290C_net ),
            .ce(),
            .sr(N__26041));
    defparam \uu2.bitmap_RNIIOM81_66_LC_5_6_0 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIIOM81_66_LC_5_6_0 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIIOM81_66_LC_5_6_0 .LUT_INIT=16'b0001000111001111;
    LogicCell40 \uu2.bitmap_RNIIOM81_66_LC_5_6_0  (
            .in0(N__13735),
            .in1(N__19436),
            .in2(N__14980),
            .in3(N__16769),
            .lcout(),
            .ltout(\uu2.bitmap_pmux_25_am_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNIM7D32_69_LC_5_6_1 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIM7D32_69_LC_5_6_1 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIM7D32_69_LC_5_6_1 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \uu2.bitmap_RNIM7D32_69_LC_5_6_1  (
            .in0(N__19437),
            .in1(N__13744),
            .in2(N__13747),
            .in3(N__14965),
            .lcout(\uu2.bitmap_RNIM7D32Z0Z_69 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_197_LC_5_6_2 .C_ON=1'b0;
    defparam \uu2.bitmap_197_LC_5_6_2 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_197_LC_5_6_2 .LUT_INIT=16'b1010101010101110;
    LogicCell40 \uu2.bitmap_197_LC_5_6_2  (
            .in0(N__19884),
            .in1(N__15060),
            .in2(N__17071),
            .in3(N__16846),
            .lcout(\uu2.bitmapZ0Z_197 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_197C_net ),
            .ce(),
            .sr(N__26039));
    defparam \uu2.bitmap_66_LC_5_6_3 .C_ON=1'b0;
    defparam \uu2.bitmap_66_LC_5_6_3 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_66_LC_5_6_3 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \uu2.bitmap_66_LC_5_6_3  (
            .in0(N__15059),
            .in1(N__19885),
            .in2(_gnd_net_),
            .in3(N__16894),
            .lcout(\uu2.bitmapZ0Z_66 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_197C_net ),
            .ce(),
            .sr(N__26039));
    defparam \uu2.bitmap_RNI2JA82_212_LC_5_6_4 .C_ON=1'b0;
    defparam \uu2.bitmap_RNI2JA82_212_LC_5_6_4 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNI2JA82_212_LC_5_6_4 .LUT_INIT=16'b0011001110111000;
    LogicCell40 \uu2.bitmap_RNI2JA82_212_LC_5_6_4  (
            .in0(N__16699),
            .in1(N__14659),
            .in2(N__16669),
            .in3(N__16770),
            .lcout(),
            .ltout(\uu2.bitmap_RNI2JA82Z0Z_212_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_nesr_RNIEE9K5_3_LC_5_6_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_RNIEE9K5_3_LC_5_6_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_nesr_RNIEE9K5_3_LC_5_6_5 .LUT_INIT=16'b0010001101100111;
    LogicCell40 \uu2.w_addr_displaying_nesr_RNIEE9K5_3_LC_5_6_5  (
            .in0(N__13725),
            .in1(N__16267),
            .in2(N__13729),
            .in3(N__13768),
            .lcout(),
            .ltout(\uu2.bitmap_pmux_27_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNI9MSLA_69_LC_5_6_6 .C_ON=1'b0;
    defparam \uu2.bitmap_RNI9MSLA_69_LC_5_6_6 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNI9MSLA_69_LC_5_6_6 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \uu2.bitmap_RNI9MSLA_69_LC_5_6_6  (
            .in0(N__13726),
            .in1(N__13714),
            .in2(N__13708),
            .in3(N__19369),
            .lcout(\uu2.N_407 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment3.segmentUQ_0_5_LC_5_7_0 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment3.segmentUQ_0_5_LC_5_7_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment3.segmentUQ_0_5_LC_5_7_0 .LUT_INIT=16'b0000110110000100;
    LogicCell40 \Lab_UT.bcd2segment3.segmentUQ_0_5_LC_5_7_0  (
            .in0(N__14763),
            .in1(N__14840),
            .in2(N__14811),
            .in3(N__14720),
            .lcout(),
            .ltout(\Lab_UT.segmentUQ_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_72_LC_5_7_1 .C_ON=1'b0;
    defparam \uu2.bitmap_72_LC_5_7_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_72_LC_5_7_1 .LUT_INIT=16'b1111111100001100;
    LogicCell40 \uu2.bitmap_72_LC_5_7_1  (
            .in0(_gnd_net_),
            .in1(N__15109),
            .in2(N__13798),
            .in3(N__19881),
            .lcout(\uu2.bitmapZ0Z_72 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_72C_net ),
            .ce(),
            .sr(N__26038));
    defparam \Lab_UT.bcd2segment3.segment_1_6_LC_5_7_2 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment3.segment_1_6_LC_5_7_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment3.segment_1_6_LC_5_7_2 .LUT_INIT=16'b1111111111011010;
    LogicCell40 \Lab_UT.bcd2segment3.segment_1_6_LC_5_7_2  (
            .in0(N__14762),
            .in1(N__14839),
            .in2(N__14810),
            .in3(N__14719),
            .lcout(\Lab_UT.segment_1_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment3.segmentUQ_i_a4_1_6_LC_5_7_3 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment3.segmentUQ_i_a4_1_6_LC_5_7_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment3.segmentUQ_i_a4_1_6_LC_5_7_3 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \Lab_UT.bcd2segment3.segmentUQ_i_a4_1_6_LC_5_7_3  (
            .in0(N__14842),
            .in1(N__14796),
            .in2(N__14728),
            .in3(N__14761),
            .lcout(),
            .ltout(\Lab_UT.N_65_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_168_LC_5_7_4 .C_ON=1'b0;
    defparam \uu2.bitmap_168_LC_5_7_4 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_168_LC_5_7_4 .LUT_INIT=16'b1010111010101010;
    LogicCell40 \uu2.bitmap_168_LC_5_7_4  (
            .in0(N__19879),
            .in1(N__15110),
            .in2(N__13795),
            .in3(N__13792),
            .lcout(\uu2.bitmapZ0Z_168 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_72C_net ),
            .ce(),
            .sr(N__26038));
    defparam \Lab_UT.bcd2segment3.segmentUQ_i_a3_4_LC_5_7_5 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment3.segmentUQ_i_a3_4_LC_5_7_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment3.segmentUQ_i_a3_4_LC_5_7_5 .LUT_INIT=16'b0000001100001010;
    LogicCell40 \Lab_UT.bcd2segment3.segmentUQ_i_a3_4_LC_5_7_5  (
            .in0(N__14841),
            .in1(N__14803),
            .in2(N__14727),
            .in3(N__14764),
            .lcout(),
            .ltout(\Lab_UT.N_76_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_200_LC_5_7_6 .C_ON=1'b0;
    defparam \uu2.bitmap_200_LC_5_7_6 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_200_LC_5_7_6 .LUT_INIT=16'b1010101010101110;
    LogicCell40 \uu2.bitmap_200_LC_5_7_6  (
            .in0(N__19880),
            .in1(N__15111),
            .in2(N__13786),
            .in3(N__13870),
            .lcout(\uu2.bitmapZ0Z_200 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_72C_net ),
            .ce(),
            .sr(N__26038));
    defparam \uu2.bitmap_RNIOS152_72_LC_5_7_7 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIOS152_72_LC_5_7_7 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIOS152_72_LC_5_7_7 .LUT_INIT=16'b0011000011101110;
    LogicCell40 \uu2.bitmap_RNIOS152_72_LC_5_7_7  (
            .in0(N__13783),
            .in1(N__19438),
            .in2(N__13777),
            .in3(N__14677),
            .lcout(\uu2.bitmap_RNIOS152Z0Z_72 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.dicLdAMtens_LC_5_8_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.dicLdAMtens_LC_5_8_0 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.dictrl.dicLdAMtens_LC_5_8_0 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \Lab_UT.dictrl.dicLdAMtens_LC_5_8_0  (
            .in0(N__20107),
            .in1(N__13921),
            .in2(N__13939),
            .in3(N__17599),
            .lcout(\Lab_UT.dictrl.dicLdAMtensZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29408),
            .ce(),
            .sr(N__13900));
    defparam \Lab_UT.didp.Mones_alarm.q_RNIN5N11_0_LC_5_8_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mones_alarm.q_RNIN5N11_0_LC_5_8_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Mones_alarm.q_RNIN5N11_0_LC_5_8_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Lab_UT.didp.Mones_alarm.q_RNIN5N11_0_LC_5_8_1  (
            .in0(N__29992),
            .in1(N__22765),
            .in2(_gnd_net_),
            .in3(N__19681),
            .lcout(\Lab_UT.Mone_at_0 ),
            .ltout(\Lab_UT.Mone_at_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment3.segmentUQ_i_a3_0_4_LC_5_8_2 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment3.segmentUQ_i_a3_0_4_LC_5_8_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment3.segmentUQ_i_a3_0_4_LC_5_8_2 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \Lab_UT.bcd2segment3.segmentUQ_i_a3_0_4_LC_5_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13873),
            .in3(N__14795),
            .lcout(\Lab_UT.N_77_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Mones_alarm.q_RNITBN11_3_LC_5_8_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mones_alarm.q_RNITBN11_3_LC_5_8_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Mones_alarm.q_RNITBN11_3_LC_5_8_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Lab_UT.didp.Mones_alarm.q_RNITBN11_3_LC_5_8_3  (
            .in0(N__28251),
            .in1(N__22693),
            .in2(_gnd_net_),
            .in3(N__19684),
            .lcout(\Lab_UT.Mone_at_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Mones_alarm.q_RNIP7N11_1_LC_5_8_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mones_alarm.q_RNIP7N11_1_LC_5_8_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Mones_alarm.q_RNIP7N11_1_LC_5_8_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.didp.Mones_alarm.q_RNIP7N11_1_LC_5_8_4  (
            .in0(N__19682),
            .in1(N__30082),
            .in2(_gnd_net_),
            .in3(N__25780),
            .lcout(\Lab_UT.Mone_at_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Mones_alarm.q_RNIR9N11_2_LC_5_8_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mones_alarm.q_RNIR9N11_2_LC_5_8_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Mones_alarm.q_RNIR9N11_2_LC_5_8_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Lab_UT.didp.Mones_alarm.q_RNIR9N11_2_LC_5_8_5  (
            .in0(N__28296),
            .in1(N__22738),
            .in2(_gnd_net_),
            .in3(N__19683),
            .lcout(\Lab_UT.Mone_at_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Mones_subtractor.q_RNIVQVP_2_LC_5_8_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mones_subtractor.q_RNIVQVP_2_LC_5_8_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Mones_subtractor.q_RNIVQVP_2_LC_5_8_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Lab_UT.didp.Mones_subtractor.q_RNIVQVP_2_LC_5_8_6  (
            .in0(N__29773),
            .in1(N__28297),
            .in2(_gnd_net_),
            .in3(N__26886),
            .lcout(\Lab_UT.didp.q_RNIVQVP_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__m22_LC_5_9_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__m22_LC_5_9_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__m22_LC_5_9_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__m22_LC_5_9_0  (
            .in0(N__23812),
            .in1(N__23976),
            .in2(_gnd_net_),
            .in3(N__15192),
            .lcout(\Lab_UT.dictrl.N_23 ),
            .ltout(\Lab_UT.dictrl.N_23_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_RNIGHD18_1_LC_5_9_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_RNIGHD18_1_LC_5_9_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_RNIGHD18_1_LC_5_9_1 .LUT_INIT=16'b0101111100001010;
    LogicCell40 \Lab_UT.dictrl.nextState_RNIGHD18_1_LC_5_9_1  (
            .in0(N__18007),
            .in1(_gnd_net_),
            .in2(N__13837),
            .in3(N__13829),
            .lcout(\Lab_UT.dictrl.nextState_RNIGHD18Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_RNIKSEU7_0_LC_5_9_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_RNIKSEU7_0_LC_5_9_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_RNIKSEU7_0_LC_5_9_2 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \Lab_UT.dictrl.currState_2_RNIKSEU7_0_LC_5_9_2  (
            .in0(N__27783),
            .in1(N__21218),
            .in2(N__15142),
            .in3(N__13804),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_12_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_RNIV4IAN_1_LC_5_9_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_RNIV4IAN_1_LC_5_9_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_RNIV4IAN_1_LC_5_9_3 .LUT_INIT=16'b1010001010000000;
    LogicCell40 \Lab_UT.dictrl.currState_2_RNIV4IAN_1_LC_5_9_3  (
            .in0(N__20188),
            .in1(N__17920),
            .in2(N__13951),
            .in3(N__17221),
            .lcout(\Lab_UT.dictrl.g0_i_a4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_RNI2P2A_2_LC_5_9_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_RNI2P2A_2_LC_5_9_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_RNI2P2A_2_LC_5_9_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Lab_UT.dictrl.currState_2_RNI2P2A_2_LC_5_9_4  (
            .in0(_gnd_net_),
            .in1(N__24964),
            .in2(_gnd_net_),
            .in3(N__23388),
            .lcout(\Lab_UT.dictrl.currState_2_RNI2P2AZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_RNI6ITB_0_2_LC_5_9_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_RNI6ITB_0_2_LC_5_9_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_RNI6ITB_0_2_LC_5_9_5 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \Lab_UT.dictrl.currState_2_RNI6ITB_0_2_LC_5_9_5  (
            .in0(N__23389),
            .in1(_gnd_net_),
            .in2(N__25009),
            .in3(N__26148),
            .lcout(\Lab_UT.dictrl.G_28_0_a5_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.dicLdAMtens_RNIDTLN4_LC_5_9_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.dicLdAMtens_RNIDTLN4_LC_5_9_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.dicLdAMtens_RNIDTLN4_LC_5_9_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \Lab_UT.dictrl.dicLdAMtens_RNIDTLN4_LC_5_9_6  (
            .in0(N__13938),
            .in1(N__13920),
            .in2(_gnd_net_),
            .in3(N__20106),
            .lcout(\Lab_UT.ld_enable_AMtens ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__m17_LC_5_9_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__m17_LC_5_9_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__m17_LC_5_9_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__m17_LC_5_9_7  (
            .in0(N__20938),
            .in1(N__27782),
            .in2(_gnd_net_),
            .in3(N__27292),
            .lcout(\Lab_UT.dictrl.N_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_0_ret_10_LC_5_10_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_10_LC_5_10_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.currState_0_ret_10_LC_5_10_0 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_10_LC_5_10_0  (
            .in0(N__14034),
            .in1(N__18009),
            .in2(N__15575),
            .in3(N__21044),
            .lcout(\Lab_UT.dictrl.r_dicLdMtens16_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29394),
            .ce(),
            .sr(N__26063));
    defparam \Lab_UT.dictrl.currState_0_ret_17_LC_5_10_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_17_LC_5_10_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.currState_0_ret_17_LC_5_10_1 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_17_LC_5_10_1  (
            .in0(N__21043),
            .in1(N__15568),
            .in2(N__18047),
            .in3(N__14035),
            .lcout(\Lab_UT.dictrl.r_dicLdMtens17_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29394),
            .ce(),
            .sr(N__26063));
    defparam \Lab_UT.dictrl.r_enable1_RNO_0_LC_5_10_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.r_enable1_RNO_0_LC_5_10_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.r_enable1_RNO_0_LC_5_10_2 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \Lab_UT.dictrl.r_enable1_RNO_0_LC_5_10_2  (
            .in0(N__15199),
            .in1(N__13909),
            .in2(_gnd_net_),
            .in3(N__17919),
            .lcout(\Lab_UT.dictrl.un1_currState_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_RNO_8_1_LC_5_10_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_RNO_8_1_LC_5_10_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_RNO_8_1_LC_5_10_3 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \Lab_UT.dictrl.nextState_RNO_8_1_LC_5_10_3  (
            .in0(N__23447),
            .in1(N__24578),
            .in2(_gnd_net_),
            .in3(N__21536),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_10_0_N_4L6_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_RNO_3_1_LC_5_10_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_RNO_3_1_LC_5_10_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_RNO_3_1_LC_5_10_4 .LUT_INIT=16'b0000000001110000;
    LogicCell40 \Lab_UT.dictrl.nextState_RNO_3_1_LC_5_10_4  (
            .in0(N__17526),
            .in1(N__15434),
            .in2(N__13903),
            .in3(N__21042),
            .lcout(\Lab_UT.dictrl.nextState_RNO_3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.r_enable4_RNO_0_LC_5_10_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.r_enable4_RNO_0_LC_5_10_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.r_enable4_RNO_0_LC_5_10_5 .LUT_INIT=16'b1010100000000000;
    LogicCell40 \Lab_UT.dictrl.r_enable4_RNO_0_LC_5_10_5  (
            .in0(N__17918),
            .in1(N__14059),
            .in2(N__14053),
            .in3(N__24863),
            .lcout(\Lab_UT.dictrl.un1_currState_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__m33_LC_5_10_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__m33_LC_5_10_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__m33_LC_5_10_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__m33_LC_5_10_6  (
            .in0(N__24862),
            .in1(N__17917),
            .in2(_gnd_net_),
            .in3(N__15181),
            .lcout(\Lab_UT.dictrl.N_34 ),
            .ltout(\Lab_UT.dictrl.N_34_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_RNIL8B7M_1_LC_5_10_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_RNIL8B7M_1_LC_5_10_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_RNIL8B7M_1_LC_5_10_7 .LUT_INIT=16'b1100111011011111;
    LogicCell40 \Lab_UT.dictrl.currState_2_RNIL8B7M_1_LC_5_10_7  (
            .in0(N__18008),
            .in1(N__24577),
            .in2(N__14038),
            .in3(N__14033),
            .lcout(\Lab_UT.dictrl.N_8ctr ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__m15_bm_LC_5_11_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__m15_bm_LC_5_11_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__m15_bm_LC_5_11_1 .LUT_INIT=16'b1101110110001101;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__m15_bm_LC_5_11_1  (
            .in0(N__17905),
            .in1(N__15211),
            .in2(N__24861),
            .in3(N__14160),
            .lcout(),
            .ltout(\Lab_UT.dictrl.m15_bm_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_0_LC_5_11_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_0_LC_5_11_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.nextState_0_LC_5_11_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \Lab_UT.dictrl.nextState_0_LC_5_11_2  (
            .in0(_gnd_net_),
            .in1(N__14113),
            .in2(N__14011),
            .in3(N__25011),
            .lcout(\Lab_UT.dictrl.nextState_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29390),
            .ce(N__15517),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_RNI1KKK6_0_LC_5_11_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_RNI1KKK6_0_LC_5_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_RNI1KKK6_0_LC_5_11_3 .LUT_INIT=16'b1111110001110100;
    LogicCell40 \Lab_UT.dictrl.nextState_RNI1KKK6_0_LC_5_11_3  (
            .in0(N__24815),
            .in1(N__18042),
            .in2(N__14007),
            .in3(N__13987),
            .lcout(\Lab_UT.dictrl.N_1609_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_3_LC_5_11_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_3_LC_5_11_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.nextState_3_LC_5_11_4 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \Lab_UT.dictrl.nextState_3_LC_5_11_4  (
            .in0(N__13975),
            .in1(N__17906),
            .in2(N__25046),
            .in3(N__23785),
            .lcout(\Lab_UT.dictrl.nextState_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29390),
            .ce(N__15517),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_ret_5_RNO_0_LC_5_11_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_ret_5_RNO_0_LC_5_11_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_ret_5_RNO_0_LC_5_11_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \Lab_UT.dictrl.currState_ret_5_RNO_0_LC_5_11_5  (
            .in0(N__23784),
            .in1(N__18084),
            .in2(_gnd_net_),
            .in3(N__23446),
            .lcout(\Lab_UT.dictrl.currState_ret_5_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_RNI1O2A_0_1_LC_5_11_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_RNI1O2A_0_1_LC_5_11_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_RNI1O2A_0_1_LC_5_11_6 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \Lab_UT.dictrl.currState_2_RNI1O2A_0_1_LC_5_11_6  (
            .in0(N__23445),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17904),
            .lcout(\Lab_UT.dictrl.currState_2_RNI1O2A_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_RNI6ITB_2_LC_5_11_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_RNI6ITB_2_LC_5_11_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_RNI6ITB_2_LC_5_11_7 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \Lab_UT.dictrl.currState_2_RNI6ITB_2_LC_5_11_7  (
            .in0(N__25010),
            .in1(N__23444),
            .in2(_gnd_net_),
            .in3(N__26147),
            .lcout(\Lab_UT.dictrl.N_23_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_16_LC_5_12_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_16_LC_5_12_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_16_LC_5_12_0 .LUT_INIT=16'b1101110111110000;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__g0_16_LC_5_12_0  (
            .in0(N__27701),
            .in1(N__21715),
            .in2(N__20398),
            .in3(N__14194),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_14_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_RNI71NQI_1_LC_5_12_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_RNI71NQI_1_LC_5_12_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_RNI71NQI_1_LC_5_12_1 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \Lab_UT.dictrl.currState_2_RNI71NQI_1_LC_5_12_1  (
            .in0(N__18062),
            .in1(N__17912),
            .in2(N__14188),
            .in3(N__14185),
            .lcout(\Lab_UT.dictrl.N_1607_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_8_LC_5_12_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_8_LC_5_12_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_8_LC_5_12_2 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__g0_8_LC_5_12_2  (
            .in0(N__20388),
            .in1(N__14175),
            .in2(_gnd_net_),
            .in3(N__14156),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_9_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_11_LC_5_12_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_11_LC_5_12_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_11_LC_5_12_3 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__g0_11_LC_5_12_3  (
            .in0(_gnd_net_),
            .in1(N__17913),
            .in2(N__14140),
            .in3(N__14131),
            .lcout(\Lab_UT.dictrl.N_10_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_6_LC_5_12_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_6_LC_5_12_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_6_LC_5_12_4 .LUT_INIT=16'b1111011100001111;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__g0_6_LC_5_12_4  (
            .in0(N__27700),
            .in1(N__14137),
            .in2(N__20397),
            .in3(N__20295),
            .lcout(\Lab_UT.dictrl.N_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__m15_am_LC_5_12_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__m15_am_LC_5_12_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__m15_am_LC_5_12_5 .LUT_INIT=16'b0111011101000100;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__m15_am_LC_5_12_5  (
            .in0(N__14125),
            .in1(N__17914),
            .in2(_gnd_net_),
            .in3(N__20283),
            .lcout(\Lab_UT.dictrl.m15_am ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_0_rep2_RNIQAFK3_LC_5_12_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_0_rep2_RNIQAFK3_LC_5_12_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_0_rep2_RNIQAFK3_LC_5_12_6 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \Lab_UT.dictrl.currState_2_0_rep2_RNIQAFK3_LC_5_12_6  (
            .in0(N__21286),
            .in1(N__18375),
            .in2(N__20939),
            .in3(N__25492),
            .lcout(\Lab_UT.dictrl.N_20_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_0_rep1_LC_5_12_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_0_rep1_LC_5_12_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.currState_2_0_rep1_LC_5_12_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Lab_UT.dictrl.currState_2_0_rep1_LC_5_12_7  (
            .in0(_gnd_net_),
            .in1(N__21071),
            .in2(_gnd_net_),
            .in3(N__24705),
            .lcout(\Lab_UT.dictrl.currState_0_rep1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29384),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.decoder.de_cr_1_0_LC_5_13_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.decoder.de_cr_1_0_LC_5_13_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.decoder.de_cr_1_0_LC_5_13_0 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \Lab_UT.dictrl.decoder.de_cr_1_0_LC_5_13_0  (
            .in0(N__15669),
            .in1(N__15681),
            .in2(_gnd_net_),
            .in3(N__14230),
            .lcout(\Lab_UT.dictrl.de_cr_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_fast_es_RNIAJ1G_3_LC_5_13_1 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_fast_es_RNIAJ1G_3_LC_5_13_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_fast_es_RNIAJ1G_3_LC_5_13_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \buart.Z_rx.bitcount_fast_es_RNIAJ1G_3_LC_5_13_1  (
            .in0(N__15673),
            .in1(N__17694),
            .in2(N__15685),
            .in3(N__15795),
            .lcout(),
            .ltout(\buart.Z_rx.bitcount_fast_es_RNIAJ1GZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_RNIK0OS_0_LC_5_13_2 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNIK0OS_0_LC_5_13_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNIK0OS_0_LC_5_13_2 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \buart.Z_rx.bitcount_es_RNIK0OS_0_LC_5_13_2  (
            .in0(N__15844),
            .in1(_gnd_net_),
            .in2(N__14275),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_rdy),
            .ltout(bu_rx_data_rdy_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_fast_RNIC98T_0_LC_5_13_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_fast_RNIC98T_0_LC_5_13_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_fast_RNIC98T_0_LC_5_13_3 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \Lab_UT.dictrl.currState_2_fast_RNIC98T_0_LC_5_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14272),
            .in3(N__14509),
            .lcout(\Lab_UT.dictrl.N_5_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__g1_0_LC_5_13_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g1_0_LC_5_13_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g1_0_LC_5_13_4 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__g1_0_LC_5_13_4  (
            .in0(N__24357),
            .in1(N__28979),
            .in2(_gnd_net_),
            .in3(N__24414),
            .lcout(\Lab_UT.dictrl.g1_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.decoder.g0_3_1_LC_5_13_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.decoder.g0_3_1_LC_5_13_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.decoder.g0_3_1_LC_5_13_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.dictrl.decoder.g0_3_1_LC_5_13_5  (
            .in0(N__28978),
            .in1(N__28606),
            .in2(_gnd_net_),
            .in3(N__24358),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_1_1_LC_5_13_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_1_1_LC_5_13_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_1_1_LC_5_13_6 .LUT_INIT=16'b0100110011001100;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__g0_1_1_LC_5_13_6  (
            .in0(N__24207),
            .in1(N__21246),
            .in2(N__14242),
            .in3(N__27712),
            .lcout(\Lab_UT.dictrl.g0_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_fast_0_LC_5_13_7 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_0_LC_5_13_7 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_fast_0_LC_5_13_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_fast_0_LC_5_13_7  (
            .in0(N__28812),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_fast_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29381),
            .ce(N__25429),
            .sr(N__26091));
    defparam \Lab_UT.dictrl.decoder.de_num_1_2_LC_5_14_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.decoder.de_num_1_2_LC_5_14_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.decoder.de_num_1_2_LC_5_14_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \Lab_UT.dictrl.decoder.de_num_1_2_LC_5_14_0  (
            .in0(N__14328),
            .in1(N__14304),
            .in2(N__14362),
            .in3(N__14313),
            .lcout(\Lab_UT.dictrl.de_num_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.decoder.g0_0_LC_5_14_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.decoder.g0_0_LC_5_14_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.decoder.g0_0_LC_5_14_1 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \Lab_UT.dictrl.decoder.g0_0_LC_5_14_1  (
            .in0(N__21895),
            .in1(N__17617),
            .in2(N__15496),
            .in3(N__14361),
            .lcout(),
            .ltout(\Lab_UT.dictrl.decoder.g0_5_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.decoder.g0_LC_5_14_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.decoder.g0_LC_5_14_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.decoder.g0_LC_5_14_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.decoder.g0_LC_5_14_2  (
            .in0(N__14338),
            .in1(N__14320),
            .in2(N__14350),
            .in3(N__17649),
            .lcout(\Lab_UT.dictrl.de_cr_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.decoder.g0_3_LC_5_14_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.decoder.g0_3_LC_5_14_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.decoder.g0_3_LC_5_14_3 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \Lab_UT.dictrl.decoder.g0_3_LC_5_14_3  (
            .in0(N__14314),
            .in1(N__20839),
            .in2(N__15843),
            .in3(N__15796),
            .lcout(\Lab_UT.dictrl.decoder.g0_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.decoder.g0_4_LC_5_14_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.decoder.g0_4_LC_5_14_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.decoder.g0_4_LC_5_14_4 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \Lab_UT.dictrl.decoder.g0_4_LC_5_14_4  (
            .in0(N__14329),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14305),
            .lcout(\Lab_UT.dictrl.decoder.g0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_fast_4_LC_5_14_5 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_4_LC_5_14_5 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_fast_4_LC_5_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_fast_4_LC_5_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24417),
            .lcout(bu_rx_data_fast_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29376),
            .ce(N__25426),
            .sr(N__26094));
    defparam \buart.Z_rx.shifter_fast_5_LC_5_14_6 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_5_LC_5_14_6 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_fast_5_LC_5_14_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_fast_5_LC_5_14_6  (
            .in0(N__24271),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_fast_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29376),
            .ce(N__25426),
            .sr(N__26094));
    defparam \buart.Z_rx.shifter_5_LC_5_14_7 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_5_LC_5_14_7 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_5_LC_5_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_5_LC_5_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24270),
            .lcout(bu_rx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29376),
            .ce(N__25426),
            .sr(N__26094));
    defparam \buart.Z_rx.hh_RNIJ3K62_0_LC_5_15_0 .C_ON=1'b0;
    defparam \buart.Z_rx.hh_RNIJ3K62_0_LC_5_15_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.hh_RNIJ3K62_0_LC_5_15_0 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \buart.Z_rx.hh_RNIJ3K62_0_LC_5_15_0  (
            .in0(N__15636),
            .in1(_gnd_net_),
            .in2(N__14296),
            .in3(N__21872),
            .lcout(\buart.Z_rx.startbit ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.decoder.g0_9_LC_5_15_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.decoder.g0_9_LC_5_15_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.decoder.g0_9_LC_5_15_1 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \Lab_UT.dictrl.decoder.g0_9_LC_5_15_1  (
            .in0(N__21764),
            .in1(N__21935),
            .in2(N__21995),
            .in3(N__17698),
            .lcout(),
            .ltout(\Lab_UT.dictrl.decoder.g0Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.decoder.g0_2_LC_5_15_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.decoder.g0_2_LC_5_15_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.decoder.g0_2_LC_5_15_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.decoder.g0_2_LC_5_15_2  (
            .in0(N__15658),
            .in1(N__14443),
            .in2(N__14512),
            .in3(N__18171),
            .lcout(\Lab_UT.dictrl.de_littleA_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__g1_4_1_LC_5_15_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g1_4_1_LC_5_15_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g1_4_1_LC_5_15_3 .LUT_INIT=16'b0101111111111111;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__g1_4_1_LC_5_15_3  (
            .in0(N__21986),
            .in1(_gnd_net_),
            .in2(N__14508),
            .in3(N__21696),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g1_4_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__g1_4_LC_5_15_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g1_4_LC_5_15_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g1_4_LC_5_15_4 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__g1_4_LC_5_15_4  (
            .in0(N__24440),
            .in1(N__21765),
            .in2(N__14467),
            .in3(N__24356),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_10_LC_5_15_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_10_LC_5_15_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_10_LC_5_15_5 .LUT_INIT=16'b1011100010111011;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__g0_10_LC_5_15_5  (
            .in0(N__24003),
            .in1(N__14464),
            .in2(N__14458),
            .in3(N__27725),
            .lcout(\Lab_UT.dictrl.N_17_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.decoder.g0_7_LC_5_15_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.decoder.g0_7_LC_5_15_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.decoder.g0_7_LC_5_15_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \Lab_UT.dictrl.decoder.g0_7_LC_5_15_6  (
            .in0(N__21394),
            .in1(N__25260),
            .in2(_gnd_net_),
            .in3(N__21697),
            .lcout(\Lab_UT.dictrl.decoder.g0_5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__m7_sx_LC_5_15_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__m7_sx_LC_5_15_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__m7_sx_LC_5_15_7 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__m7_sx_LC_5_15_7  (
            .in0(N__21763),
            .in1(N__21695),
            .in2(N__24012),
            .in3(N__21393),
            .lcout(\Lab_UT.dictrl.m7_sx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_0_LC_5_16_3 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_0_LC_5_16_3 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_0_LC_5_16_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_0_LC_5_16_3  (
            .in0(_gnd_net_),
            .in1(N__15922),
            .in2(_gnd_net_),
            .in3(N__14414),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29371),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_RNI3O55_3_LC_5_16_5 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI3O55_3_LC_5_16_5 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI3O55_3_LC_5_16_5 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_RNI3O55_3_LC_5_16_5  (
            .in0(N__14427),
            .in1(N__14413),
            .in2(_gnd_net_),
            .in3(N__14395),
            .lcout(\buart.Z_rx.ser_clk ),
            .ltout(\buart.Z_rx.ser_clk_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_4_LC_5_16_6 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_4_LC_5_16_6 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_4_LC_5_16_6 .LUT_INIT=16'b0000000100000100;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_4_LC_5_16_6  (
            .in0(N__15921),
            .in1(N__14389),
            .in2(N__14383),
            .in3(N__14379),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29371),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_RNIGD8S2_1_LC_5_16_7 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNIGD8S2_1_LC_5_16_7 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNIGD8S2_1_LC_5_16_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \buart.Z_rx.bitcount_es_RNIGD8S2_1_LC_5_16_7  (
            .in0(N__15637),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27729),
            .lcout(\buart.Z_rx.N_27_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_0_LC_6_3_0 .C_ON=1'b0;
    defparam \resetGen.reset_count_0_LC_6_3_0 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_0_LC_6_3_0 .LUT_INIT=16'b0000000010011001;
    LogicCell40 \resetGen.reset_count_0_LC_6_3_0  (
            .in0(N__19172),
            .in1(N__19218),
            .in2(_gnd_net_),
            .in3(N__20433),
            .lcout(\resetGen.reset_countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29437),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_RNO_0_4_LC_6_3_1 .C_ON=1'b0;
    defparam \resetGen.reset_count_RNO_0_4_LC_6_3_1 .SEQ_MODE=4'b0000;
    defparam \resetGen.reset_count_RNO_0_4_LC_6_3_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \resetGen.reset_count_RNO_0_4_LC_6_3_1  (
            .in0(_gnd_net_),
            .in1(N__18937),
            .in2(_gnd_net_),
            .in3(N__19144),
            .lcout(),
            .ltout(\resetGen.reset_count_2_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_4_LC_6_3_2 .C_ON=1'b0;
    defparam \resetGen.reset_count_4_LC_6_3_2 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_4_LC_6_3_2 .LUT_INIT=16'b0000000011101100;
    LogicCell40 \resetGen.reset_count_4_LC_6_3_2  (
            .in0(N__19204),
            .in1(N__19171),
            .in2(N__14566),
            .in3(N__20434),
            .lcout(\resetGen.reset_countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29437),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_1_LC_6_3_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_1_LC_6_3_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_1_LC_6_3_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_1_LC_6_3_3  (
            .in0(N__19035),
            .in1(N__18771),
            .in2(_gnd_net_),
            .in3(N__14917),
            .lcout(\uu2.mem0.w_addr_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_3_LC_6_3_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_3_LC_6_3_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_3_LC_6_3_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_3_LC_6_3_4  (
            .in0(N__18772),
            .in1(N__22460),
            .in2(_gnd_net_),
            .in3(N__16505),
            .lcout(\uu2.mem0.w_addr_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_6__un426_ci_3_LC_6_3_5 .C_ON=1'b0;
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_6__un426_ci_3_LC_6_3_5 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_6__un426_ci_3_LC_6_3_5 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \uu2.vbuf_w_addr_user.counter_gen_label_6__un426_ci_3_LC_6_3_5  (
            .in0(N__22461),
            .in1(_gnd_net_),
            .in2(N__22492),
            .in3(_gnd_net_),
            .lcout(\uu2.un426_ci_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_4_LC_6_3_6 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_4_LC_6_3_6 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_4_LC_6_3_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_4_LC_6_3_6  (
            .in0(N__18773),
            .in1(N__22488),
            .in2(_gnd_net_),
            .in3(N__16543),
            .lcout(\uu2.mem0.w_addr_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_5_LC_6_3_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_5_LC_6_3_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_5_LC_6_3_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_5_LC_6_3_7  (
            .in0(N__22351),
            .in1(N__16446),
            .in2(_gnd_net_),
            .in3(N__18774),
            .lcout(\uu2.mem0.w_addr_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIGEPH1_4_LC_6_4_0 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIGEPH1_4_LC_6_4_0 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIGEPH1_4_LC_6_4_0 .LUT_INIT=16'b0101110010000000;
    LogicCell40 \uu2.w_addr_displaying_RNIGEPH1_4_LC_6_4_0  (
            .in0(N__16256),
            .in1(N__16504),
            .in2(N__16121),
            .in3(N__14909),
            .lcout(\uu2.bitmap_pmux_sn_N_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNI6RO21_162_LC_6_4_1 .C_ON=1'b0;
    defparam \uu2.bitmap_RNI6RO21_162_LC_6_4_1 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNI6RO21_162_LC_6_4_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \uu2.bitmap_RNI6RO21_162_LC_6_4_1  (
            .in0(N__14620),
            .in1(N__16253),
            .in2(_gnd_net_),
            .in3(N__14938),
            .lcout(),
            .ltout(\uu2.N_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNIELSJ2_111_LC_6_4_2 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIELSJ2_111_LC_6_4_2 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIELSJ2_111_LC_6_4_2 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \uu2.bitmap_RNIELSJ2_111_LC_6_4_2  (
            .in0(_gnd_net_),
            .in1(N__14596),
            .in2(N__14611),
            .in3(N__14602),
            .lcout(\uu2.bitmap_RNIELSJ2Z0Z_111 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIM0T61_2_LC_6_4_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIM0T61_2_LC_6_4_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIM0T61_2_LC_6_4_3 .LUT_INIT=16'b1010101000010001;
    LogicCell40 \uu2.w_addr_displaying_RNIM0T61_2_LC_6_4_3  (
            .in0(N__14907),
            .in1(N__16254),
            .in2(_gnd_net_),
            .in3(N__16103),
            .lcout(\uu2.bitmap_pmux_sn_N_54_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_111_LC_6_4_4 .C_ON=1'b0;
    defparam \uu2.bitmap_111_LC_6_4_4 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_111_LC_6_4_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.bitmap_111_LC_6_4_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26800),
            .lcout(\uu2.bitmapZ0Z_111 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_111C_net ),
            .ce(),
            .sr(N__26046));
    defparam \uu2.w_addr_displaying_RNI8NSO_4_LC_6_4_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI8NSO_4_LC_6_4_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI8NSO_4_LC_6_4_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.w_addr_displaying_RNI8NSO_4_LC_6_4_5  (
            .in0(_gnd_net_),
            .in1(N__16498),
            .in2(_gnd_net_),
            .in3(N__16104),
            .lcout(\uu2.bitmap_pmux_sn_N_33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI8NSO_2_LC_6_4_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI8NSO_2_LC_6_4_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI8NSO_2_LC_6_4_6 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \uu2.w_addr_displaying_RNI8NSO_2_LC_6_4_6  (
            .in0(N__16255),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14908),
            .lcout(\uu2.N_39 ),
            .ltout(\uu2.N_39_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_w_addr_displaying.result_1_0_o2_4_LC_6_4_7 .C_ON=1'b0;
    defparam \uu2.vbuf_w_addr_displaying.result_1_0_o2_4_LC_6_4_7 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_w_addr_displaying.result_1_0_o2_4_LC_6_4_7 .LUT_INIT=16'b1111001111111111;
    LogicCell40 \uu2.vbuf_w_addr_displaying.result_1_0_o2_4_LC_6_4_7  (
            .in0(_gnd_net_),
            .in1(N__19496),
            .in2(N__14569),
            .in3(N__16108),
            .lcout(\uu2.N_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_nesr_3_LC_6_5_0 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_3_LC_6_5_0 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_nesr_3_LC_6_5_0 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.w_addr_displaying_nesr_3_LC_6_5_0  (
            .in0(N__16120),
            .in1(N__14906),
            .in2(N__19497),
            .in3(N__16271),
            .lcout(\uu2.w_addr_displayingZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_nesr_3C_net ),
            .ce(N__16303),
            .sr(N__26044));
    defparam \uu2.w_addr_displaying_nesr_1_LC_6_5_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_1_LC_6_5_1 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_nesr_1_LC_6_5_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.w_addr_displaying_nesr_1_LC_6_5_1  (
            .in0(_gnd_net_),
            .in1(N__19483),
            .in2(_gnd_net_),
            .in3(N__16119),
            .lcout(\uu2.w_addr_displayingZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_nesr_3C_net ),
            .ce(N__16303),
            .sr(N__26044));
    defparam \uu2.w_addr_displaying_nesr_7_LC_6_5_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_7_LC_6_5_2 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_nesr_7_LC_6_5_2 .LUT_INIT=16'b1010100110101010;
    LogicCell40 \uu2.w_addr_displaying_nesr_7_LC_6_5_2  (
            .in0(N__16778),
            .in1(N__16461),
            .in2(N__16374),
            .in3(N__16441),
            .lcout(\uu2.w_addr_displayingZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_nesr_3C_net ),
            .ce(N__16303),
            .sr(N__26044));
    defparam \uu2.w_addr_displaying_ness_6_LC_6_5_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_ness_6_LC_6_5_3 .SEQ_MODE=4'b1001;
    defparam \uu2.w_addr_displaying_ness_6_LC_6_5_3 .LUT_INIT=16'b1010101011010101;
    LogicCell40 \uu2.w_addr_displaying_ness_6_LC_6_5_3  (
            .in0(N__16440),
            .in1(N__16777),
            .in2(N__16639),
            .in3(N__14671),
            .lcout(\uu2.w_addr_displayingZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_nesr_3C_net ),
            .ce(N__16303),
            .sr(N__26044));
    defparam CONSTANT_ONE_LUT4_LC_6_5_4.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_6_5_4.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_6_5_4.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_6_5_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNI35M31_84_LC_6_6_0 .C_ON=1'b0;
    defparam \uu2.bitmap_RNI35M31_84_LC_6_6_0 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNI35M31_84_LC_6_6_0 .LUT_INIT=16'b0010010100101111;
    LogicCell40 \uu2.bitmap_RNI35M31_84_LC_6_6_0  (
            .in0(N__16757),
            .in1(N__14653),
            .in2(N__19459),
            .in3(N__16900),
            .lcout(\uu2.bitmap_pmux_24_am_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_87_LC_6_6_1 .C_ON=1'b0;
    defparam \uu2.bitmap_87_LC_6_6_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_87_LC_6_6_1 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \uu2.bitmap_87_LC_6_6_1  (
            .in0(N__19882),
            .in1(N__16294),
            .in2(_gnd_net_),
            .in3(N__20170),
            .lcout(\uu2.bitmapZ0Z_87 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_87C_net ),
            .ce(),
            .sr(N__26042));
    defparam \uu2.bitmap_314_LC_6_6_2 .C_ON=1'b0;
    defparam \uu2.bitmap_314_LC_6_6_2 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_314_LC_6_6_2 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \uu2.bitmap_314_LC_6_6_2  (
            .in0(N__19543),
            .in1(N__19883),
            .in2(_gnd_net_),
            .in3(N__19096),
            .lcout(\uu2.bitmapZ0Z_314 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_87C_net ),
            .ce(),
            .sr(N__26042));
    defparam \uu2.bitmap_RNIVKR41_180_LC_6_6_3 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIVKR41_180_LC_6_6_3 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIVKR41_180_LC_6_6_3 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \uu2.bitmap_RNIVKR41_180_LC_6_6_3  (
            .in0(_gnd_net_),
            .in1(N__16678),
            .in2(N__16272),
            .in3(N__14640),
            .lcout(),
            .ltout(\uu2.N_386_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_nesr_RNI1JET2_7_LC_6_6_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_RNI1JET2_7_LC_6_6_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_nesr_RNI1JET2_7_LC_6_6_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \uu2.w_addr_displaying_nesr_RNI1JET2_7_LC_6_6_4  (
            .in0(N__16756),
            .in1(N__16250),
            .in2(N__14647),
            .in3(N__16558),
            .lcout(),
            .ltout(\uu2.w_addr_displaying_nesr_RNI1JET2Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNIMAS54_314_LC_6_6_5 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIMAS54_314_LC_6_6_5 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIMAS54_314_LC_6_6_5 .LUT_INIT=16'b0000110100101111;
    LogicCell40 \uu2.bitmap_RNIMAS54_314_LC_6_6_5  (
            .in0(N__16252),
            .in1(N__16110),
            .in2(N__14644),
            .in3(N__14641),
            .lcout(\uu2.bitmap_pmux_23_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIAGTK1_2_LC_6_6_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIAGTK1_2_LC_6_6_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIAGTK1_2_LC_6_6_6 .LUT_INIT=16'b0000011100000110;
    LogicCell40 \uu2.w_addr_displaying_RNIAGTK1_2_LC_6_6_6  (
            .in0(N__14898),
            .in1(N__16109),
            .in2(N__16779),
            .in3(N__16251),
            .lcout(\uu2.bitmap_pmux_sn_N_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_2_LC_6_6_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_2_LC_6_6_7 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_2_LC_6_6_7 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu2.w_addr_displaying_2_LC_6_6_7  (
            .in0(N__19473),
            .in1(N__14899),
            .in2(N__16336),
            .in3(N__16111),
            .lcout(\uu2.w_addr_displayingZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_87C_net ),
            .ce(),
            .sr(N__26042));
    defparam \Lab_UT.didp.Mones_alarm.q_RNI83T64_1_1_LC_6_7_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mones_alarm.q_RNI83T64_1_1_LC_6_7_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Mones_alarm.q_RNI83T64_1_1_LC_6_7_0 .LUT_INIT=16'b0000100010010010;
    LogicCell40 \Lab_UT.didp.Mones_alarm.q_RNI83T64_1_1_LC_6_7_0  (
            .in0(N__14835),
            .in1(N__14804),
            .in2(N__14765),
            .in3(N__14715),
            .lcout(\Lab_UT.L3_segment3_0_i_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Mones_alarm.q_RNI83T64_1_LC_6_7_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mones_alarm.q_RNI83T64_1_LC_6_7_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Mones_alarm.q_RNI83T64_1_LC_6_7_1 .LUT_INIT=16'b0110011011011011;
    LogicCell40 \Lab_UT.didp.Mones_alarm.q_RNI83T64_1_LC_6_7_1  (
            .in0(N__14716),
            .in1(N__14754),
            .in2(N__14812),
            .in3(N__14836),
            .lcout(\Lab_UT.L3_segment3_0_i_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Mones_alarm.q_RNI83T64_0_1_LC_6_7_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mones_alarm.q_RNI83T64_0_1_LC_6_7_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Mones_alarm.q_RNI83T64_0_1_LC_6_7_2 .LUT_INIT=16'b0011111010111111;
    LogicCell40 \Lab_UT.didp.Mones_alarm.q_RNI83T64_0_1_LC_6_7_2  (
            .in0(N__14837),
            .in1(N__14808),
            .in2(N__14766),
            .in3(N__14717),
            .lcout(),
            .ltout(\Lab_UT.L3_segment3_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_203_LC_6_7_3 .C_ON=1'b0;
    defparam \uu2.bitmap_203_LC_6_7_3 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_203_LC_6_7_3 .LUT_INIT=16'b0000000011000000;
    LogicCell40 \uu2.bitmap_203_LC_6_7_3  (
            .in0(_gnd_net_),
            .in1(N__15107),
            .in2(N__14845),
            .in3(N__19893),
            .lcout(\uu2.bitmapZ0Z_203 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_203C_net ),
            .ce(),
            .sr(N__26040));
    defparam \Lab_UT.didp.Mones_alarm.q_RNI83T64_2_1_LC_6_7_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mones_alarm.q_RNI83T64_2_1_LC_6_7_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Mones_alarm.q_RNI83T64_2_1_LC_6_7_4 .LUT_INIT=16'b0010011110011111;
    LogicCell40 \Lab_UT.didp.Mones_alarm.q_RNI83T64_2_1_LC_6_7_4  (
            .in0(N__14838),
            .in1(N__14809),
            .in2(N__14767),
            .in3(N__14718),
            .lcout(),
            .ltout(\Lab_UT.L3_segment3_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_75_LC_6_7_5 .C_ON=1'b0;
    defparam \uu2.bitmap_75_LC_6_7_5 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_75_LC_6_7_5 .LUT_INIT=16'b0000000011000000;
    LogicCell40 \uu2.bitmap_75_LC_6_7_5  (
            .in0(_gnd_net_),
            .in1(N__15108),
            .in2(N__14692),
            .in3(N__19894),
            .lcout(\uu2.bitmapZ0Z_75 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_203C_net ),
            .ce(),
            .sr(N__26040));
    defparam \uu2.bitmap_RNI99H91_75_LC_6_7_6 .C_ON=1'b0;
    defparam \uu2.bitmap_RNI99H91_75_LC_6_7_6 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNI99H91_75_LC_6_7_6 .LUT_INIT=16'b0011000001011111;
    LogicCell40 \uu2.bitmap_RNI99H91_75_LC_6_7_6  (
            .in0(N__14689),
            .in1(N__14683),
            .in2(N__19458),
            .in3(N__16780),
            .lcout(\uu2.bitmap_pmux_24_bm_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_0_LC_6_7_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_0_LC_6_7_7 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_0_LC_6_7_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \uu2.w_addr_displaying_0_LC_6_7_7  (
            .in0(N__16332),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19425),
            .lcout(\uu2.w_addr_displayingZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_203C_net ),
            .ce(),
            .sr(N__26040));
    defparam \Lab_UT.bcd2segment4.segmentUQ_i_a3_4_LC_6_8_0 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment4.segmentUQ_i_a3_4_LC_6_8_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment4.segmentUQ_i_a3_4_LC_6_8_0 .LUT_INIT=16'b0000000000101110;
    LogicCell40 \Lab_UT.bcd2segment4.segmentUQ_i_a3_4_LC_6_8_0  (
            .in0(N__17041),
            .in1(N__19604),
            .in2(N__17001),
            .in3(N__16940),
            .lcout(),
            .ltout(\Lab_UT.N_76_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_194_LC_6_8_1 .C_ON=1'b0;
    defparam \uu2.bitmap_194_LC_6_8_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_194_LC_6_8_1 .LUT_INIT=16'b1111111100000100;
    LogicCell40 \uu2.bitmap_194_LC_6_8_1  (
            .in0(N__16948),
            .in1(N__15055),
            .in2(N__14983),
            .in3(N__19896),
            .lcout(\uu2.bitmapZ0Z_194 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_194C_net ),
            .ce(),
            .sr(N__26037));
    defparam \Lab_UT.didp.Mtens_alarm.q_RNIGGJ64_2_LC_6_8_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mtens_alarm.q_RNIGGJ64_2_LC_6_8_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Mtens_alarm.q_RNIGGJ64_2_LC_6_8_2 .LUT_INIT=16'b0010000010000110;
    LogicCell40 \Lab_UT.didp.Mtens_alarm.q_RNIGGJ64_2_LC_6_8_2  (
            .in0(N__17040),
            .in1(N__19603),
            .in2(N__17000),
            .in3(N__16939),
            .lcout(\Lab_UT.L3_segment4_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Mtens_alarm.q_RNIGGJ64_0_2_LC_6_8_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mtens_alarm.q_RNIGGJ64_0_2_LC_6_8_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Mtens_alarm.q_RNIGGJ64_0_2_LC_6_8_3 .LUT_INIT=16'b0110011100011111;
    LogicCell40 \Lab_UT.didp.Mtens_alarm.q_RNIGGJ64_0_2_LC_6_8_3  (
            .in0(N__16941),
            .in1(N__16994),
            .in2(N__19609),
            .in3(N__17042),
            .lcout(),
            .ltout(\Lab_UT.L3_segment4_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_69_LC_6_8_4 .C_ON=1'b0;
    defparam \uu2.bitmap_69_LC_6_8_4 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_69_LC_6_8_4 .LUT_INIT=16'b0000000011000000;
    LogicCell40 \uu2.bitmap_69_LC_6_8_4  (
            .in0(_gnd_net_),
            .in1(N__15039),
            .in2(N__14968),
            .in3(N__19820),
            .lcout(\uu2.bitmapZ0Z_69 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_194C_net ),
            .ce(),
            .sr(N__26037));
    defparam \uu2.bitmap_34_LC_6_8_5 .C_ON=1'b0;
    defparam \uu2.bitmap_34_LC_6_8_5 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_34_LC_6_8_5 .LUT_INIT=16'b0000000000001010;
    LogicCell40 \uu2.bitmap_34_LC_6_8_5  (
            .in0(N__15038),
            .in1(_gnd_net_),
            .in2(N__19875),
            .in3(N__14956),
            .lcout(\uu2.bitmapZ0Z_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_194C_net ),
            .ce(),
            .sr(N__26037));
    defparam \Lab_UT.bcd2segment4.segment_1_6_LC_6_8_6 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment4.segment_1_6_LC_6_8_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment4.segment_1_6_LC_6_8_6 .LUT_INIT=16'b1111111110111100;
    LogicCell40 \Lab_UT.bcd2segment4.segment_1_6_LC_6_8_6  (
            .in0(N__17043),
            .in1(N__19608),
            .in2(N__17002),
            .in3(N__16942),
            .lcout(),
            .ltout(\Lab_UT.segment_1_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_162_LC_6_8_7 .C_ON=1'b0;
    defparam \uu2.bitmap_162_LC_6_8_7 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_162_LC_6_8_7 .LUT_INIT=16'b1100110011101100;
    LogicCell40 \uu2.bitmap_162_LC_6_8_7  (
            .in0(N__15040),
            .in1(N__19895),
            .in2(N__14941),
            .in3(N__16882),
            .lcout(\uu2.bitmapZ0Z_162 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_194C_net ),
            .ce(),
            .sr(N__26037));
    defparam \Lab_UT.dictrl.nextState_RNI6VQ05_2_LC_6_9_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_RNI6VQ05_2_LC_6_9_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_RNI6VQ05_2_LC_6_9_0 .LUT_INIT=16'b1100110010100000;
    LogicCell40 \Lab_UT.dictrl.nextState_RNI6VQ05_2_LC_6_9_0  (
            .in0(N__18130),
            .in1(N__15537),
            .in2(N__20857),
            .in3(N__23436),
            .lcout(\Lab_UT.dictrl.N_1614_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_0_ret_21_RNIUL8L_LC_6_9_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_21_RNIUL8L_LC_6_9_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_0_ret_21_RNIUL8L_LC_6_9_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_21_RNIUL8L_LC_6_9_1  (
            .in0(N__18013),
            .in1(N__23813),
            .in2(_gnd_net_),
            .in3(N__24006),
            .lcout(\Lab_UT.dictrl.N_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.r_enable1_LC_6_9_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.r_enable1_LC_6_9_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.r_enable1_LC_6_9_2 .LUT_INIT=16'b1100111111001010;
    LogicCell40 \Lab_UT.dictrl.r_enable1_LC_6_9_2  (
            .in0(N__15133),
            .in1(N__15127),
            .in2(N__23457),
            .in3(N__20200),
            .lcout(\Lab_UT.dictrl.r_enableZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29393),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.r_enable1_RNI7DR61_LC_6_9_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.r_enable1_RNI7DR61_LC_6_9_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.r_enable1_RNI7DR61_LC_6_9_3 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \Lab_UT.dictrl.r_enable1_RNI7DR61_LC_6_9_3  (
            .in0(N__15126),
            .in1(N__24168),
            .in2(N__23176),
            .in3(N__23654),
            .lcout(\Lab_UT.dictrl.enableSeg1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.r_enable3_RNI9DR61_LC_6_9_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.r_enable3_RNI9DR61_LC_6_9_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.r_enable3_RNI9DR61_LC_6_9_4 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \Lab_UT.dictrl.r_enable3_RNI9DR61_LC_6_9_4  (
            .in0(N__23655),
            .in1(N__15072),
            .in2(N__24176),
            .in3(N__23174),
            .lcout(\Lab_UT.dictrl.enableSeg3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.r_enable3_LC_6_9_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.r_enable3_LC_6_9_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.r_enable3_LC_6_9_5 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \Lab_UT.dictrl.r_enable3_LC_6_9_5  (
            .in0(N__23437),
            .in1(N__19695),
            .in2(N__15076),
            .in3(N__21307),
            .lcout(\Lab_UT.dictrl.r_enableZ0Z3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29393),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.r_enable4_RNIADR61_LC_6_9_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.r_enable4_RNIADR61_LC_6_9_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.r_enable4_RNIADR61_LC_6_9_6 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \Lab_UT.dictrl.r_enable4_RNIADR61_LC_6_9_6  (
            .in0(N__23656),
            .in1(N__15000),
            .in2(N__24177),
            .in3(N__23175),
            .lcout(\Lab_UT.dictrl.enableSeg4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.r_enable4_LC_6_9_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.r_enable4_LC_6_9_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.r_enable4_LC_6_9_7 .LUT_INIT=16'b1010000010110001;
    LogicCell40 \Lab_UT.dictrl.r_enable4_LC_6_9_7  (
            .in0(N__23438),
            .in1(N__19696),
            .in2(N__15004),
            .in3(N__15013),
            .lcout(\Lab_UT.dictrl.r_enableZ0Z4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29393),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_RNI19TAN_1_LC_6_10_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_RNI19TAN_1_LC_6_10_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_RNI19TAN_1_LC_6_10_0 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \Lab_UT.dictrl.currState_2_RNI19TAN_1_LC_6_10_0  (
            .in0(N__14992),
            .in1(N__17911),
            .in2(_gnd_net_),
            .in3(N__17230),
            .lcout(\Lab_UT.dictrl.g1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_RNI421C4_0_LC_6_10_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_RNI421C4_0_LC_6_10_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_RNI421C4_0_LC_6_10_1 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \Lab_UT.dictrl.currState_2_RNI421C4_0_LC_6_10_1  (
            .in0(N__27285),
            .in1(N__21250),
            .in2(N__27810),
            .in3(N__17442),
            .lcout(\Lab_UT.dictrl.N_17_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_19_LC_6_10_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_19_LC_6_10_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_19_LC_6_10_2 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__g0_19_LC_6_10_2  (
            .in0(N__17629),
            .in1(N__27777),
            .in2(N__21264),
            .in3(N__27284),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_36_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_RNIBR9BG_1_LC_6_10_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_RNIBR9BG_1_LC_6_10_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_RNIBR9BG_1_LC_6_10_3 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \Lab_UT.dictrl.currState_2_RNIBR9BG_1_LC_6_10_3  (
            .in0(_gnd_net_),
            .in1(N__17443),
            .in2(N__15205),
            .in3(N__17452),
            .lcout(\Lab_UT.dictrl.nextStateZ0Z_3 ),
            .ltout(\Lab_UT.dictrl.nextStateZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_0_ret_26_LC_6_10_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_26_LC_6_10_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.currState_0_ret_26_LC_6_10_4 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_26_LC_6_10_4  (
            .in0(_gnd_net_),
            .in1(N__24682),
            .in2(N__15202),
            .in3(N__21072),
            .lcout(\Lab_UT.dictrl.r_dicLdMtens21_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29388),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_0_ret_25_LC_6_10_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_25_LC_6_10_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.currState_0_ret_25_LC_6_10_5 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_25_LC_6_10_5  (
            .in0(N__17546),
            .in1(N__15474),
            .in2(N__17356),
            .in3(N__15385),
            .lcout(\Lab_UT.dictrl.r_dicLdMtens22_i_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29388),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_0_ret_27_LC_6_10_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_27_LC_6_10_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.currState_0_ret_27_LC_6_10_6 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_27_LC_6_10_6  (
            .in0(N__15475),
            .in1(N__17355),
            .in2(N__17335),
            .in3(N__17547),
            .lcout(\Lab_UT.dictrl.r_dicLdMtens20_i_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29388),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__m32_LC_6_10_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__m32_LC_6_10_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__m32_LC_6_10_7 .LUT_INIT=16'b0010000001110101;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__m32_LC_6_10_7  (
            .in0(N__23816),
            .in1(N__24481),
            .in2(N__21265),
            .in3(N__15193),
            .lcout(\Lab_UT.dictrl.N_33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_RNIDED951_2_LC_6_11_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_RNIDED951_2_LC_6_11_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_RNIDED951_2_LC_6_11_0 .LUT_INIT=16'b1100100011001101;
    LogicCell40 \Lab_UT.dictrl.currState_2_RNIDED951_2_LC_6_11_0  (
            .in0(N__23453),
            .in1(N__15175),
            .in2(N__25047),
            .in3(N__15169),
            .lcout(\Lab_UT.dictrl.nextStateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_RNID73K33_1_LC_6_11_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_RNID73K33_1_LC_6_11_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_RNID73K33_1_LC_6_11_1 .LUT_INIT=16'b1111011101111111;
    LogicCell40 \Lab_UT.dictrl.currState_2_RNID73K33_1_LC_6_11_1  (
            .in0(N__21035),
            .in1(N__15163),
            .in2(N__21609),
            .in3(N__20751),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_0_ret_29_RNIOSJNC6_LC_6_11_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_29_RNIOSJNC6_LC_6_11_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_0_ret_29_RNIOSJNC6_LC_6_11_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_29_RNIOSJNC6_LC_6_11_2  (
            .in0(N__23454),
            .in1(N__24677),
            .in2(N__15286),
            .in3(N__17128),
            .lcout(\Lab_UT.dictrl.g0_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_RNO_9_1_LC_6_11_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_RNO_9_1_LC_6_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_RNO_9_1_LC_6_11_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \Lab_UT.dictrl.nextState_RNO_9_1_LC_6_11_3  (
            .in0(N__24678),
            .in1(N__23455),
            .in2(_gnd_net_),
            .in3(N__20668),
            .lcout(),
            .ltout(\Lab_UT.dictrl.nextState_RNO_9Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_RNO_4_1_LC_6_11_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_RNO_4_1_LC_6_11_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_RNO_4_1_LC_6_11_4 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \Lab_UT.dictrl.nextState_RNO_4_1_LC_6_11_4  (
            .in0(N__15279),
            .in1(N__15244),
            .in2(N__15283),
            .in3(N__17122),
            .lcout(),
            .ltout(\Lab_UT.dictrl.nextState_RNO_4Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_RNO_1_1_LC_6_11_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_RNO_1_1_LC_6_11_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_RNO_1_1_LC_6_11_5 .LUT_INIT=16'b0000000001110000;
    LogicCell40 \Lab_UT.dictrl.nextState_RNO_1_1_LC_6_11_5  (
            .in0(N__15280),
            .in1(N__15238),
            .in2(N__15262),
            .in3(N__15259),
            .lcout(\Lab_UT.dictrl.g0_i_o4_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_RNO_11_1_LC_6_11_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_RNO_11_1_LC_6_11_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_RNO_11_1_LC_6_11_6 .LUT_INIT=16'b1100000011001111;
    LogicCell40 \Lab_UT.dictrl.nextState_RNO_11_1_LC_6_11_6  (
            .in0(_gnd_net_),
            .in1(N__21568),
            .in2(N__20795),
            .in3(N__21036),
            .lcout(\Lab_UT.dictrl.N_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_RNO_5_1_LC_6_11_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_RNO_5_1_LC_6_11_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_RNO_5_1_LC_6_11_7 .LUT_INIT=16'b0001000000110000;
    LogicCell40 \Lab_UT.dictrl.nextState_RNO_5_1_LC_6_11_7  (
            .in0(N__17532),
            .in1(N__20755),
            .in2(N__21610),
            .in3(N__15484),
            .lcout(\Lab_UT.dictrl.N_18_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_23_LC_6_12_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_23_LC_6_12_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_23_LC_6_12_0 .LUT_INIT=16'b0111001011111010;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__g0_23_LC_6_12_0  (
            .in0(N__21259),
            .in1(N__27710),
            .in2(N__18343),
            .in3(N__27299),
            .lcout(\Lab_UT.dictrl.N_13_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__g1_LC_6_12_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g1_LC_6_12_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g1_LC_6_12_1 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__g1_LC_6_12_1  (
            .in0(N__23831),
            .in1(N__24309),
            .in2(N__15232),
            .in3(N__28602),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g1_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_22_LC_6_12_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_22_LC_6_12_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_22_LC_6_12_2 .LUT_INIT=16'b1110010011101110;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__g0_22_LC_6_12_2  (
            .in0(N__15223),
            .in1(N__23832),
            .in2(N__15214),
            .in3(N__27711),
            .lcout(\Lab_UT.dictrl.N_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_0_ret_28_RNO_0_LC_6_12_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_28_RNO_0_LC_6_12_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_0_ret_28_RNO_0_LC_6_12_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_28_RNO_0_LC_6_12_3  (
            .in0(N__17351),
            .in1(N__17553),
            .in2(N__17331),
            .in3(N__15481),
            .lcout(),
            .ltout(\Lab_UT.dictrl.r_dicLdMtens20_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_0_ret_28_LC_6_12_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_28_LC_6_12_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.currState_0_ret_28_LC_6_12_4 .LUT_INIT=16'b0000010000001100;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_28_LC_6_12_4  (
            .in0(N__15409),
            .in1(N__17488),
            .in2(N__15487),
            .in3(N__15358),
            .lcout(\Lab_UT.dictrl.r_Sone_init17_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29379),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_RNIFGT042_0_LC_6_12_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_RNIFGT042_0_LC_6_12_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_RNIFGT042_0_LC_6_12_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.dictrl.currState_2_RNIFGT042_0_LC_6_12_5  (
            .in0(_gnd_net_),
            .in1(N__17552),
            .in2(_gnd_net_),
            .in3(N__15480),
            .lcout(\Lab_UT.dictrl.r_dicLdMtens22_2_reti ),
            .ltout(\Lab_UT.dictrl.r_dicLdMtens22_2_reti_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_0_ret_29_RNIDFRSEE_LC_6_12_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_29_RNIDFRSEE_LC_6_12_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_0_ret_29_RNIDFRSEE_LC_6_12_6 .LUT_INIT=16'b0001010100000000;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_29_RNIDFRSEE_LC_6_12_6  (
            .in0(N__15403),
            .in1(N__15357),
            .in2(N__15394),
            .in3(N__15391),
            .lcout(\Lab_UT.dictrl.currState_0_ret_29_RNIDFRSEEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_0_ret_21_RNIPJM6D1_LC_6_12_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_21_RNIPJM6D1_LC_6_12_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_0_ret_21_RNIPJM6D1_LC_6_12_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_21_RNIPJM6D1_LC_6_12_7  (
            .in0(N__17350),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15384),
            .lcout(\Lab_UT.dictrl.r_dicLdMtens22_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__m27_LC_6_13_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__m27_LC_6_13_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__m27_LC_6_13_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__m27_LC_6_13_0  (
            .in0(N__15297),
            .in1(N__21267),
            .in2(_gnd_net_),
            .in3(N__24874),
            .lcout(\Lab_UT.dictrl.N_41_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_RNIN9NP3_7_LC_6_13_1 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_RNIN9NP3_7_LC_6_13_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.shifter_RNIN9NP3_7_LC_6_13_1 .LUT_INIT=16'b1011111111111111;
    LogicCell40 \buart.Z_rx.shifter_RNIN9NP3_7_LC_6_13_1  (
            .in0(N__25397),
            .in1(N__21290),
            .in2(N__18376),
            .in3(N__25478),
            .lcout(N_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__m29_LC_6_13_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__m29_LC_6_13_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__m29_LC_6_13_2 .LUT_INIT=16'b0010011110101111;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__m29_LC_6_13_2  (
            .in0(N__23798),
            .in1(N__17099),
            .in2(N__15337),
            .in3(N__21266),
            .lcout(\Lab_UT.dictrl.N_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.decoder.de_littleA_LC_6_13_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.decoder.de_littleA_LC_6_13_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.decoder.de_littleA_LC_6_13_3 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \Lab_UT.dictrl.decoder.de_littleA_LC_6_13_3  (
            .in0(N__25398),
            .in1(N__17473),
            .in2(N__24208),
            .in3(N__21291),
            .lcout(\Lab_UT.dictrl.de_littleA ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.decoder.de_cr_1_LC_6_13_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.decoder.de_cr_1_LC_6_13_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.decoder.de_cr_1_LC_6_13_4 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \Lab_UT.dictrl.decoder.de_cr_1_LC_6_13_4  (
            .in0(N__18224),
            .in1(N__18179),
            .in2(_gnd_net_),
            .in3(N__17650),
            .lcout(Lab_UT_dictrl_decoder_de_cr_1),
            .ltout(Lab_UT_dictrl_decoder_de_cr_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.decoder.de_cr_LC_6_13_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.decoder.de_cr_LC_6_13_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.decoder.de_cr_LC_6_13_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \Lab_UT.dictrl.decoder.de_cr_LC_6_13_5  (
            .in0(N__18371),
            .in1(N__25394),
            .in2(N__15598),
            .in3(N__25477),
            .lcout(\Lab_UT.dictrl.de_cr ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__m30_LC_6_13_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__m30_LC_6_13_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__m30_LC_6_13_6 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__m30_LC_6_13_6  (
            .in0(N__17928),
            .in1(N__15595),
            .in2(_gnd_net_),
            .in3(N__15589),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_2_LC_6_13_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_2_LC_6_13_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.nextState_2_LC_6_13_7 .LUT_INIT=16'b1100110000001111;
    LogicCell40 \Lab_UT.dictrl.nextState_2_LC_6_13_7  (
            .in0(_gnd_net_),
            .in1(N__15582),
            .in2(N__15544),
            .in3(N__25040),
            .lcout(\Lab_UT.dictrl.nextState_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29374),
            .ce(N__15513),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_fast_es_2_LC_6_14_0 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_fast_es_2_LC_6_14_0 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_fast_es_2_LC_6_14_0 .LUT_INIT=16'b0010011101110010;
    LogicCell40 \buart.Z_rx.bitcount_fast_es_2_LC_6_14_0  (
            .in0(N__15977),
            .in1(N__15931),
            .in2(N__15745),
            .in3(N__18236),
            .lcout(buart__rx_bitcount_fast_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29372),
            .ce(N__15870),
            .sr(N__26095));
    defparam \buart.Z_rx.bitcount_es_2_LC_6_14_1 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_2_LC_6_14_1 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_es_2_LC_6_14_1 .LUT_INIT=16'b0001110100101110;
    LogicCell40 \buart.Z_rx.bitcount_es_2_LC_6_14_1  (
            .in0(N__18235),
            .in1(N__15974),
            .in2(N__15941),
            .in3(N__15740),
            .lcout(buart__rx_bitcount_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29372),
            .ce(N__15870),
            .sr(N__26095));
    defparam \buart.Z_rx.bitcount_2_rep1_es_LC_6_14_2 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_2_rep1_es_LC_6_14_2 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_2_rep1_es_LC_6_14_2 .LUT_INIT=16'b0010011101110010;
    LogicCell40 \buart.Z_rx.bitcount_2_rep1_es_LC_6_14_2  (
            .in0(N__15972),
            .in1(N__15928),
            .in2(N__15744),
            .in3(N__18234),
            .lcout(buart__rx_bitcount_2_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29372),
            .ce(N__15870),
            .sr(N__26095));
    defparam \buart.Z_rx.bitcount_es_1_LC_6_14_3 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_1_LC_6_14_3 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_es_1_LC_6_14_3 .LUT_INIT=16'b0100011101110100;
    LogicCell40 \buart.Z_rx.bitcount_es_1_LC_6_14_3  (
            .in0(N__15927),
            .in1(N__15973),
            .in2(N__15760),
            .in3(N__15803),
            .lcout(buart__rx_bitcount_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29372),
            .ce(N__15870),
            .sr(N__26095));
    defparam \buart.Z_rx.bitcount_es_4_LC_6_14_4 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_4_LC_6_14_4 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_es_4_LC_6_14_4 .LUT_INIT=16'b0010011101110010;
    LogicCell40 \buart.Z_rx.bitcount_es_4_LC_6_14_4  (
            .in0(N__15976),
            .in1(N__15930),
            .in2(N__15700),
            .in3(N__18319),
            .lcout(buart__rx_bitcount_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29372),
            .ce(N__15870),
            .sr(N__26095));
    defparam \buart.Z_rx.bitcount_fast_es_4_LC_6_14_5 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_fast_es_4_LC_6_14_5 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_fast_es_4_LC_6_14_5 .LUT_INIT=16'b0001110100101110;
    LogicCell40 \buart.Z_rx.bitcount_fast_es_4_LC_6_14_5  (
            .in0(N__18318),
            .in1(N__15979),
            .in2(N__15943),
            .in3(N__15699),
            .lcout(buart__rx_bitcount_fast_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29372),
            .ce(N__15870),
            .sr(N__26095));
    defparam \buart.Z_rx.bitcount_es_3_LC_6_14_6 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_3_LC_6_14_6 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_es_3_LC_6_14_6 .LUT_INIT=16'b0010011101110010;
    LogicCell40 \buart.Z_rx.bitcount_es_3_LC_6_14_6  (
            .in0(N__15975),
            .in1(N__15929),
            .in2(N__15721),
            .in3(N__18278),
            .lcout(buart__rx_bitcount_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29372),
            .ce(N__15870),
            .sr(N__26095));
    defparam \buart.Z_rx.bitcount_fast_es_3_LC_6_14_7 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_fast_es_3_LC_6_14_7 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_fast_es_3_LC_6_14_7 .LUT_INIT=16'b0001110100101110;
    LogicCell40 \buart.Z_rx.bitcount_fast_es_3_LC_6_14_7  (
            .in0(N__18279),
            .in1(N__15978),
            .in2(N__15942),
            .in3(N__15720),
            .lcout(buart__rx_bitcount_fast_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29372),
            .ce(N__15870),
            .sr(N__26095));
    defparam \Lab_UT.dictrl.decoder.g0_8_LC_6_15_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.decoder.g0_8_LC_6_15_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.decoder.g0_8_LC_6_15_0 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Lab_UT.dictrl.decoder.g0_8_LC_6_15_0  (
            .in0(N__18269),
            .in1(N__21837),
            .in2(N__18321),
            .in3(N__21351),
            .lcout(\Lab_UT.dictrl.decoder.g0_6_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_RNIIVPI1_1_LC_6_15_1 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNIIVPI1_1_LC_6_15_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNIIVPI1_1_LC_6_15_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \buart.Z_rx.bitcount_es_RNIIVPI1_1_LC_6_15_1  (
            .in0(N__18232),
            .in1(N__18270),
            .in2(N__15804),
            .in3(N__18317),
            .lcout(),
            .ltout(\buart.Z_rx.un1_sample_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_RNIV4M42_0_LC_6_15_2 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNIV4M42_0_LC_6_15_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNIV4M42_0_LC_6_15_2 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \buart.Z_rx.bitcount_es_RNIV4M42_0_LC_6_15_2  (
            .in0(N__15837),
            .in1(_gnd_net_),
            .in2(N__15652),
            .in3(N__15619),
            .lcout(\buart.Z_rx.sample ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_RNILRCP_0_LC_6_15_3 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNILRCP_0_LC_6_15_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNILRCP_0_LC_6_15_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \buart.Z_rx.bitcount_es_RNILRCP_0_LC_6_15_3  (
            .in0(_gnd_net_),
            .in1(N__15835),
            .in2(_gnd_net_),
            .in3(N__15793),
            .lcout(buart__rx_valid_2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_RNIOUCP_0_LC_6_15_4 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNIOUCP_0_LC_6_15_4 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNIOUCP_0_LC_6_15_4 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \buart.Z_rx.bitcount_es_RNIOUCP_0_LC_6_15_4  (
            .in0(N__15836),
            .in1(_gnd_net_),
            .in2(N__18322),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\buart.Z_rx.idle_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_RNISCGV1_1_LC_6_15_5 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNISCGV1_1_LC_6_15_5 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNISCGV1_1_LC_6_15_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \buart.Z_rx.bitcount_es_RNISCGV1_1_LC_6_15_5  (
            .in0(N__18233),
            .in1(N__18271),
            .in2(N__15640),
            .in3(N__15794),
            .lcout(\buart.Z_rx.idle ),
            .ltout(\buart.Z_rx.idle_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_fast_sbtinv_3_LC_6_15_6 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_fast_sbtinv_3_LC_6_15_6 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_fast_sbtinv_3_LC_6_15_6 .LUT_INIT=16'b1111111110101110;
    LogicCell40 \buart.Z_rx.bitcount_fast_sbtinv_3_LC_6_15_6  (
            .in0(N__15919),
            .in1(N__15620),
            .in2(N__15601),
            .in3(N__27781),
            .lcout(\buart.Z_rx.bitcounte_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_0_LC_6_15_7 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_0_LC_6_15_7 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_es_0_LC_6_15_7 .LUT_INIT=16'b0010011101110010;
    LogicCell40 \buart.Z_rx.bitcount_es_0_LC_6_15_7  (
            .in0(N__15954),
            .in1(N__15920),
            .in2(N__28356),
            .in3(N__15838),
            .lcout(buart__rx_bitcount_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29370),
            .ce(N__15871),
            .sr(N__26096));
    defparam \buart.Z_rx.bitcount_cry_c_0_LC_6_16_0 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_c_0_LC_6_16_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_c_0_LC_6_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_c_0_LC_6_16_0  (
            .in0(_gnd_net_),
            .in1(N__15842),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_16_0_),
            .carryout(\buart.Z_rx.bitcount_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_6_16_1 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_6_16_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_6_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_6_16_1  (
            .in0(_gnd_net_),
            .in1(N__15805),
            .in2(_gnd_net_),
            .in3(N__15748),
            .lcout(\buart.Z_rx.bitcount_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.bitcount_cry_0 ),
            .carryout(\buart.Z_rx.bitcount_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_6_16_2 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_6_16_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_6_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_6_16_2  (
            .in0(_gnd_net_),
            .in1(N__18238),
            .in2(_gnd_net_),
            .in3(N__15724),
            .lcout(\buart.Z_rx.bitcount_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.bitcount_cry_1 ),
            .carryout(\buart.Z_rx.bitcount_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_6_16_3 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_6_16_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_6_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_6_16_3  (
            .in0(_gnd_net_),
            .in1(N__18280),
            .in2(_gnd_net_),
            .in3(N__15706),
            .lcout(\buart.Z_rx.bitcount_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.bitcount_cry_2 ),
            .carryout(\buart.Z_rx.bitcount_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_3_THRU_LUT4_0_LC_6_16_4 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_cry_3_THRU_LUT4_0_LC_6_16_4 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_3_THRU_LUT4_0_LC_6_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_3_THRU_LUT4_0_LC_6_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15703),
            .lcout(\buart.Z_rx.bitcount_cry_3_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.decoder.g0_3_0_LC_6_16_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.decoder.g0_3_0_LC_6_16_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.decoder.g0_3_0_LC_6_16_6 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \Lab_UT.dictrl.decoder.g0_3_0_LC_6_16_6  (
            .in0(N__28974),
            .in1(N__18237),
            .in2(_gnd_net_),
            .in3(N__28601),
            .lcout(\Lab_UT.dictrl.decoder.g0_3Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.uu0.l_count_18_LC_7_1_0 .C_ON=1'b0;
    defparam \Lab_UT.uu0.l_count_18_LC_7_1_0 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.uu0.l_count_18_LC_7_1_0 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \Lab_UT.uu0.l_count_18_LC_7_1_0  (
            .in0(N__18460),
            .in1(N__22071),
            .in2(_gnd_net_),
            .in3(N__23248),
            .lcout(\Lab_UT.uu0.l_countZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29463),
            .ce(N__22174),
            .sr(N__26099));
    defparam \Lab_UT.uu0.l_count_13_LC_7_1_4 .C_ON=1'b0;
    defparam \Lab_UT.uu0.l_count_13_LC_7_1_4 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.uu0.l_count_13_LC_7_1_4 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \Lab_UT.uu0.l_count_13_LC_7_1_4  (
            .in0(N__18602),
            .in1(N__16029),
            .in2(N__15988),
            .in3(N__23247),
            .lcout(\Lab_UT.uu0.l_countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29463),
            .ce(N__22174),
            .sr(N__26099));
    defparam \Lab_UT.uu0.l_count_2_LC_7_1_6 .C_ON=1'b0;
    defparam \Lab_UT.uu0.l_count_2_LC_7_1_6 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.uu0.l_count_2_LC_7_1_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Lab_UT.uu0.l_count_2_LC_7_1_6  (
            .in0(_gnd_net_),
            .in1(N__21793),
            .in2(_gnd_net_),
            .in3(N__22241),
            .lcout(\Lab_UT.uu0.l_countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29463),
            .ce(N__22174),
            .sr(N__26099));
    defparam \Lab_UT.uu0.l_count_RNIFRMN_3_LC_7_2_0 .C_ON=1'b0;
    defparam \Lab_UT.uu0.l_count_RNIFRMN_3_LC_7_2_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.uu0.l_count_RNIFRMN_3_LC_7_2_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \Lab_UT.uu0.l_count_RNIFRMN_3_LC_7_2_0  (
            .in0(N__18450),
            .in1(N__18500),
            .in2(N__18487),
            .in3(N__22264),
            .lcout(\Lab_UT.uu0.un4_l_count_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.uu0.l_count_12_LC_7_2_1 .C_ON=1'b0;
    defparam \Lab_UT.uu0.l_count_12_LC_7_2_1 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.uu0.l_count_12_LC_7_2_1 .LUT_INIT=16'b0001001000100010;
    LogicCell40 \Lab_UT.uu0.l_count_12_LC_7_2_1  (
            .in0(N__16005),
            .in1(N__23240),
            .in2(N__18694),
            .in3(N__18604),
            .lcout(\Lab_UT.uu0.l_countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29456),
            .ce(N__22172),
            .sr(N__26098));
    defparam \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_7_2_2 .C_ON=1'b0;
    defparam \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_7_2_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_7_2_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_7_2_2  (
            .in0(N__18558),
            .in1(N__18452),
            .in2(_gnd_net_),
            .in3(N__18430),
            .lcout(),
            .ltout(\Lab_UT.uu0.un143_ci_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.uu0.l_count_11_LC_7_2_3 .C_ON=1'b0;
    defparam \Lab_UT.uu0.l_count_11_LC_7_2_3 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.uu0.l_count_11_LC_7_2_3 .LUT_INIT=16'b0001001000100010;
    LogicCell40 \Lab_UT.uu0.l_count_11_LC_7_2_3  (
            .in0(N__22560),
            .in1(N__23239),
            .in2(N__16015),
            .in3(N__18603),
            .lcout(\Lab_UT.uu0.l_countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29456),
            .ce(N__22172),
            .sr(N__26098));
    defparam \Lab_UT.uu0.l_count_9_LC_7_2_4 .C_ON=1'b0;
    defparam \Lab_UT.uu0.l_count_9_LC_7_2_4 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.uu0.l_count_9_LC_7_2_4 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \Lab_UT.uu0.l_count_9_LC_7_2_4  (
            .in0(N__18559),
            .in1(_gnd_net_),
            .in2(N__18610),
            .in3(N__18453),
            .lcout(\Lab_UT.uu0.l_countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29456),
            .ce(N__22172),
            .sr(N__26098));
    defparam \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_7_2_5 .C_ON=1'b0;
    defparam \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_7_2_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_7_2_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_7_2_5  (
            .in0(N__18451),
            .in1(N__18429),
            .in2(N__22561),
            .in3(N__18557),
            .lcout(\Lab_UT.uu0.un154_ci_9 ),
            .ltout(\Lab_UT.uu0.un154_ci_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_7_2_6 .C_ON=1'b0;
    defparam \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_7_2_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_7_2_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_7_2_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16012),
            .in3(N__16004),
            .lcout(\Lab_UT.uu0.un165_ci_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_RNI1VU6_3_LC_7_3_0 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_RNI1VU6_3_LC_7_3_0 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_nesr_RNI1VU6_3_LC_7_3_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uu2.w_addr_user_nesr_RNI1VU6_3_LC_7_3_0  (
            .in0(N__22487),
            .in1(N__18991),
            .in2(N__16155),
            .in3(N__19049),
            .lcout(\uu2.un3_w_addr_user_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_RNI7UV5_8_LC_7_3_1 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_RNI7UV5_8_LC_7_3_1 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_nesr_RNI7UV5_8_LC_7_3_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \uu2.w_addr_user_nesr_RNI7UV5_8_LC_7_3_1  (
            .in0(N__22459),
            .in1(N__16172),
            .in2(_gnd_net_),
            .in3(N__18962),
            .lcout(),
            .ltout(\uu2.un3_w_addr_user_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_RNIINVH_2_LC_7_3_2 .C_ON=1'b0;
    defparam \uu2.w_addr_user_RNIINVH_2_LC_7_3_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_RNIINVH_2_LC_7_3_2 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \uu2.w_addr_user_RNIINVH_2_LC_7_3_2  (
            .in0(N__22352),
            .in1(N__19030),
            .in2(N__16285),
            .in3(N__16282),
            .lcout(\uu2.un3_w_addr_user ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_3_LC_7_3_3 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_3_LC_7_3_3 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_nesr_3_LC_7_3_3 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu2.w_addr_user_nesr_3_LC_7_3_3  (
            .in0(N__19050),
            .in1(N__18993),
            .in2(N__19036),
            .in3(N__18963),
            .lcout(\uu2.w_addr_userZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_nesr_3C_net ),
            .ce(N__18535),
            .sr(N__22322));
    defparam \uu2.mem0.ram512X8_inst_RNO_2_LC_7_3_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_2_LC_7_3_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_2_LC_7_3_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_2_LC_7_3_4  (
            .in0(N__18992),
            .in1(N__18749),
            .in2(_gnd_net_),
            .in3(N__16276),
            .lcout(\uu2.mem0.w_addr_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_8__un448_ci_0_LC_7_3_5 .C_ON=1'b0;
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_8__un448_ci_0_LC_7_3_5 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_8__un448_ci_0_LC_7_3_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.vbuf_w_addr_user.counter_gen_label_8__un448_ci_0_LC_7_3_5  (
            .in0(_gnd_net_),
            .in1(N__22353),
            .in2(_gnd_net_),
            .in3(N__16150),
            .lcout(),
            .ltout(\uu2.vbuf_w_addr_user.un448_ci_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_8_LC_7_3_6 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_8_LC_7_3_6 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_nesr_8_LC_7_3_6 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \uu2.w_addr_user_nesr_8_LC_7_3_6  (
            .in0(N__16173),
            .in1(N__22370),
            .in2(N__16180),
            .in3(N__22399),
            .lcout(\uu2.w_addr_userZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_nesr_3C_net ),
            .ce(N__18535),
            .sr(N__22322));
    defparam \uu2.w_addr_user_nesr_7_LC_7_3_7 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_7_LC_7_3_7 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_nesr_7_LC_7_3_7 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.w_addr_user_nesr_7_LC_7_3_7  (
            .in0(N__22398),
            .in1(N__22354),
            .in2(N__22374),
            .in3(N__16151),
            .lcout(\uu2.w_addr_userZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_nesr_3C_net ),
            .ce(N__18535),
            .sr(N__22322));
    defparam \uu2.w_addr_displaying_RNIHGM43_8_LC_7_4_0 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIHGM43_8_LC_7_4_0 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIHGM43_8_LC_7_4_0 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \uu2.w_addr_displaying_RNIHGM43_8_LC_7_4_0  (
            .in0(N__16118),
            .in1(N__16388),
            .in2(N__16052),
            .in3(N__16616),
            .lcout(\uu2.N_71 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_8_LC_7_4_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_8_LC_7_4_1 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_8_LC_7_4_1 .LUT_INIT=16'b1100110011000110;
    LogicCell40 \uu2.w_addr_displaying_8_LC_7_4_1  (
            .in0(N__16331),
            .in1(N__16618),
            .in2(N__16397),
            .in3(N__16364),
            .lcout(\uu2.w_addr_displayingZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_8C_net ),
            .ce(),
            .sr(N__26049));
    defparam \uu2.w_addr_displaying_4_LC_7_4_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_4_LC_7_4_2 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_4_LC_7_4_2 .LUT_INIT=16'b1011101101000100;
    LogicCell40 \uu2.w_addr_displaying_4_LC_7_4_2  (
            .in0(N__16362),
            .in1(N__16329),
            .in2(_gnd_net_),
            .in3(N__16500),
            .lcout(\uu2.w_addr_displayingZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_8C_net ),
            .ce(),
            .sr(N__26049));
    defparam \uu2.w_addr_displaying_5_LC_7_4_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_5_LC_7_4_3 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_5_LC_7_4_3 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \uu2.w_addr_displaying_5_LC_7_4_3  (
            .in0(N__16330),
            .in1(N__16506),
            .in2(N__16544),
            .in3(N__16363),
            .lcout(\uu2.w_addr_displayingZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_8C_net ),
            .ce(),
            .sr(N__26049));
    defparam \uu2.w_addr_displaying_RNILSOL_5_LC_7_4_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNILSOL_5_LC_7_4_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNILSOL_5_LC_7_4_4 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \uu2.w_addr_displaying_RNILSOL_5_LC_7_4_4  (
            .in0(_gnd_net_),
            .in1(N__16533),
            .in2(_gnd_net_),
            .in3(N__16499),
            .lcout(\uu2.N_41 ),
            .ltout(\uu2.N_41_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_ness_RNITTSI1_6_LC_7_4_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_ness_RNITTSI1_6_LC_7_4_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_ness_RNITTSI1_6_LC_7_4_5 .LUT_INIT=16'b1111001111111111;
    LogicCell40 \uu2.w_addr_displaying_ness_RNITTSI1_6_LC_7_4_5  (
            .in0(_gnd_net_),
            .in1(N__16433),
            .in2(N__16402),
            .in3(N__16771),
            .lcout(\uu2.N_43 ),
            .ltout(\uu2.N_43_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIFCPV4_8_LC_7_4_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIFCPV4_8_LC_7_4_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIFCPV4_8_LC_7_4_6 .LUT_INIT=16'b0011011100110011;
    LogicCell40 \uu2.w_addr_displaying_RNIFCPV4_8_LC_7_4_6  (
            .in0(N__16361),
            .in1(N__18748),
            .in2(N__16339),
            .in3(N__16617),
            .lcout(\uu2.w_addr_displaying_RNIFCPV4Z0Z_8 ),
            .ltout(\uu2.w_addr_displaying_RNIFCPV4Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIJ5K15_8_LC_7_4_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIJ5K15_8_LC_7_4_7 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIJ5K15_8_LC_7_4_7 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \uu2.w_addr_displaying_RNIJ5K15_8_LC_7_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16306),
            .in3(N__26146),
            .lcout(\uu2.N_36_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Stens_alarm.q_RNI0QLC5_2_1_LC_7_5_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.Stens_alarm.q_RNI0QLC5_2_1_LC_7_5_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Stens_alarm.q_RNI0QLC5_2_1_LC_7_5_0 .LUT_INIT=16'b0001101110110111;
    LogicCell40 \Lab_UT.didp.Stens_alarm.q_RNI0QLC5_2_1_LC_7_5_0  (
            .in0(N__20044),
            .in1(N__19938),
            .in2(N__20008),
            .in3(N__20074),
            .lcout(\Lab_UT.L3_segment2_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Stens_alarm.q_RNI0QLC5_1_LC_7_5_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.Stens_alarm.q_RNI0QLC5_1_LC_7_5_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Stens_alarm.q_RNI0QLC5_1_LC_7_5_1 .LUT_INIT=16'b0101101011100111;
    LogicCell40 \Lab_UT.didp.Stens_alarm.q_RNI0QLC5_1_LC_7_5_1  (
            .in0(N__20077),
            .in1(N__20007),
            .in2(N__19951),
            .in3(N__20047),
            .lcout(),
            .ltout(\Lab_UT.L3_segment2_0_i_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_308_LC_7_5_2 .C_ON=1'b0;
    defparam \uu2.bitmap_308_LC_7_5_2 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_308_LC_7_5_2 .LUT_INIT=16'b1111101010101010;
    LogicCell40 \uu2.bitmap_308_LC_7_5_2  (
            .in0(N__19849),
            .in1(_gnd_net_),
            .in2(N__16288),
            .in3(N__20168),
            .lcout(\uu2.bitmapZ0Z_308 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_308C_net ),
            .ce(),
            .sr(N__26047));
    defparam \Lab_UT.didp.Stens_alarm.q_RNI0QLC5_0_1_LC_7_5_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.Stens_alarm.q_RNI0QLC5_0_1_LC_7_5_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Stens_alarm.q_RNI0QLC5_0_1_LC_7_5_3 .LUT_INIT=16'b0111111100111101;
    LogicCell40 \Lab_UT.didp.Stens_alarm.q_RNI0QLC5_0_1_LC_7_5_3  (
            .in0(N__20075),
            .in1(N__20005),
            .in2(N__19949),
            .in3(N__20045),
            .lcout(),
            .ltout(\Lab_UT.L3_segment2_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_215_LC_7_5_4 .C_ON=1'b0;
    defparam \uu2.bitmap_215_LC_7_5_4 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_215_LC_7_5_4 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \uu2.bitmap_215_LC_7_5_4  (
            .in0(N__19848),
            .in1(_gnd_net_),
            .in2(N__16672),
            .in3(N__20167),
            .lcout(\uu2.bitmapZ0Z_215 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_308C_net ),
            .ce(),
            .sr(N__26047));
    defparam \Lab_UT.didp.Stens_alarm.q_RNI0QLC5_1_1_LC_7_5_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.Stens_alarm.q_RNI0QLC5_1_1_LC_7_5_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Stens_alarm.q_RNI0QLC5_1_1_LC_7_5_5 .LUT_INIT=16'b0100100100010000;
    LogicCell40 \Lab_UT.didp.Stens_alarm.q_RNI0QLC5_1_1_LC_7_5_5  (
            .in0(N__20076),
            .in1(N__20006),
            .in2(N__19950),
            .in3(N__20046),
            .lcout(),
            .ltout(\Lab_UT.L3_segment2_0_i_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_52_LC_7_5_6 .C_ON=1'b0;
    defparam \uu2.bitmap_52_LC_7_5_6 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_52_LC_7_5_6 .LUT_INIT=16'b1010111110101010;
    LogicCell40 \uu2.bitmap_52_LC_7_5_6  (
            .in0(N__19850),
            .in1(_gnd_net_),
            .in2(N__16654),
            .in3(N__20169),
            .lcout(\uu2.bitmapZ0Z_52 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_308C_net ),
            .ce(),
            .sr(N__26047));
    defparam \uu2.bitmap_RNIU2IS_52_LC_7_5_7 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIU2IS_52_LC_7_5_7 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIU2IS_52_LC_7_5_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \uu2.bitmap_RNIU2IS_52_LC_7_5_7  (
            .in0(N__16651),
            .in1(N__16604),
            .in2(_gnd_net_),
            .in3(N__16564),
            .lcout(\uu2.N_158 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.segmentUQ_0_5_LC_7_6_0 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.segmentUQ_0_5_LC_7_6_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.segmentUQ_0_5_LC_7_6_0 .LUT_INIT=16'b0010100000110010;
    LogicCell40 \Lab_UT.bcd2segment1.segmentUQ_0_5_LC_7_6_0  (
            .in0(N__19358),
            .in1(N__19311),
            .in2(N__19741),
            .in3(N__19269),
            .lcout(),
            .ltout(\Lab_UT.segmentUQ_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_90_LC_7_6_1 .C_ON=1'b0;
    defparam \uu2.bitmap_90_LC_7_6_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_90_LC_7_6_1 .LUT_INIT=16'b1100111111001100;
    LogicCell40 \uu2.bitmap_90_LC_7_6_1  (
            .in0(_gnd_net_),
            .in1(N__19886),
            .in2(N__16552),
            .in3(N__19559),
            .lcout(\uu2.bitmapZ0Z_90 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_90C_net ),
            .ce(),
            .sr(N__26045));
    defparam \Lab_UT.bcd2segment1.segment_1_6_LC_7_6_2 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.segment_1_6_LC_7_6_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.segment_1_6_LC_7_6_2 .LUT_INIT=16'b1111101111111100;
    LogicCell40 \Lab_UT.bcd2segment1.segment_1_6_LC_7_6_2  (
            .in0(N__19357),
            .in1(N__19310),
            .in2(N__19740),
            .in3(N__19268),
            .lcout(\Lab_UT.segment_1_2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.segmentUQ_i_a4_1_6_LC_7_6_3 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.segmentUQ_i_a4_1_6_LC_7_6_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.segmentUQ_i_a4_1_6_LC_7_6_3 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \Lab_UT.bcd2segment1.segmentUQ_i_a4_1_6_LC_7_6_3  (
            .in0(N__19267),
            .in1(N__19737),
            .in2(N__19317),
            .in3(N__19360),
            .lcout(),
            .ltout(\Lab_UT.N_65_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_186_LC_7_6_4 .C_ON=1'b0;
    defparam \uu2.bitmap_186_LC_7_6_4 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_186_LC_7_6_4 .LUT_INIT=16'b1100111011001100;
    LogicCell40 \uu2.bitmap_186_LC_7_6_4  (
            .in0(N__19560),
            .in1(N__19855),
            .in2(N__16825),
            .in3(N__16822),
            .lcout(\uu2.bitmapZ0Z_186 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_90C_net ),
            .ce(),
            .sr(N__26045));
    defparam \Lab_UT.bcd2segment1.segmentUQ_i_a3_4_LC_7_6_5 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.segmentUQ_i_a3_4_LC_7_6_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.segmentUQ_i_a3_4_LC_7_6_5 .LUT_INIT=16'b0001001100000010;
    LogicCell40 \Lab_UT.bcd2segment1.segmentUQ_i_a3_4_LC_7_6_5  (
            .in0(N__19270),
            .in1(N__19736),
            .in2(N__19318),
            .in3(N__19359),
            .lcout(),
            .ltout(\Lab_UT.N_76_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_218_LC_7_6_6 .C_ON=1'b0;
    defparam \uu2.bitmap_218_LC_7_6_6 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_218_LC_7_6_6 .LUT_INIT=16'b1100110111001100;
    LogicCell40 \uu2.bitmap_218_LC_7_6_6  (
            .in0(N__19327),
            .in1(N__19856),
            .in2(N__16807),
            .in3(N__19564),
            .lcout(\uu2.bitmapZ0Z_218 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_90C_net ),
            .ce(),
            .sr(N__26045));
    defparam \uu2.bitmap_RNICFK91_90_LC_7_6_7 .C_ON=1'b0;
    defparam \uu2.bitmap_RNICFK91_90_LC_7_6_7 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNICFK91_90_LC_7_6_7 .LUT_INIT=16'b0001000111001111;
    LogicCell40 \uu2.bitmap_RNICFK91_90_LC_7_6_7  (
            .in0(N__16804),
            .in1(N__19435),
            .in2(N__16798),
            .in3(N__16767),
            .lcout(\uu2.bitmap_pmux_25_bm_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment2.segment_1_6_LC_7_7_0 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment2.segment_1_6_LC_7_7_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment2.segment_1_6_LC_7_7_0 .LUT_INIT=16'b1111111110111100;
    LogicCell40 \Lab_UT.bcd2segment2.segment_1_6_LC_7_7_0  (
            .in0(N__20041),
            .in1(N__19983),
            .in2(N__19948),
            .in3(N__20071),
            .lcout(\Lab_UT.segment_1_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment2.segmentUQ_i_a3_4_LC_7_7_1 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment2.segmentUQ_i_a3_4_LC_7_7_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment2.segmentUQ_i_a3_4_LC_7_7_1 .LUT_INIT=16'b0001010100000100;
    LogicCell40 \Lab_UT.bcd2segment2.segmentUQ_i_a3_4_LC_7_7_1  (
            .in0(N__20072),
            .in1(N__19937),
            .in2(N__19992),
            .in3(N__20042),
            .lcout(),
            .ltout(\Lab_UT.N_76_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_212_LC_7_7_2 .C_ON=1'b0;
    defparam \uu2.bitmap_212_LC_7_7_2 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_212_LC_7_7_2 .LUT_INIT=16'b1100110011001110;
    LogicCell40 \uu2.bitmap_212_LC_7_7_2  (
            .in0(N__20166),
            .in1(N__19878),
            .in2(N__16702),
            .in3(N__16906),
            .lcout(\uu2.bitmapZ0Z_212 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_212C_net ),
            .ce(),
            .sr(N__26043));
    defparam \Lab_UT.bcd2segment2.segmentUQ_i_a4_1_6_LC_7_7_3 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment2.segmentUQ_i_a4_1_6_LC_7_7_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment2.segmentUQ_i_a4_1_6_LC_7_7_3 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \Lab_UT.bcd2segment2.segmentUQ_i_a4_1_6_LC_7_7_3  (
            .in0(N__20073),
            .in1(N__19933),
            .in2(N__19991),
            .in3(N__20043),
            .lcout(),
            .ltout(\Lab_UT.N_65_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_180_LC_7_7_4 .C_ON=1'b0;
    defparam \uu2.bitmap_180_LC_7_7_4 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_180_LC_7_7_4 .LUT_INIT=16'b1100111011001100;
    LogicCell40 \uu2.bitmap_180_LC_7_7_4  (
            .in0(N__20165),
            .in1(N__19877),
            .in2(N__16687),
            .in3(N__16684),
            .lcout(\uu2.bitmapZ0Z_180 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_212C_net ),
            .ce(),
            .sr(N__26043));
    defparam \Lab_UT.bcd2segment2.segmentUQ_i_a3_0_4_LC_7_7_5 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment2.segmentUQ_i_a3_0_4_LC_7_7_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment2.segmentUQ_i_a3_0_4_LC_7_7_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.bcd2segment2.segmentUQ_i_a3_0_4_LC_7_7_5  (
            .in0(_gnd_net_),
            .in1(N__19979),
            .in2(_gnd_net_),
            .in3(N__20040),
            .lcout(\Lab_UT.N_77_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_84_LC_7_7_7 .C_ON=1'b0;
    defparam \uu2.bitmap_84_LC_7_7_7 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_84_LC_7_7_7 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \uu2.bitmap_84_LC_7_7_7  (
            .in0(N__19876),
            .in1(N__20164),
            .in2(_gnd_net_),
            .in3(N__19903),
            .lcout(\uu2.bitmapZ0Z_84 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_212C_net ),
            .ce(),
            .sr(N__26043));
    defparam \Lab_UT.didp.Mtens_alarm.q_RNIO8T96_3_LC_7_8_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mtens_alarm.q_RNIO8T96_3_LC_7_8_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Mtens_alarm.q_RNIO8T96_3_LC_7_8_0 .LUT_INIT=16'b0110011001101111;
    LogicCell40 \Lab_UT.didp.Mtens_alarm.q_RNIO8T96_3_LC_7_8_0  (
            .in0(N__16834),
            .in1(N__16979),
            .in2(N__17044),
            .in3(N__16857),
            .lcout(\Lab_UT.L3_segment4_0_i_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment4.segmentUQ_i_a4_1_6_LC_7_8_1 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment4.segmentUQ_i_a4_1_6_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment4.segmentUQ_i_a4_1_6_LC_7_8_1 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \Lab_UT.bcd2segment4.segmentUQ_i_a4_1_6_LC_7_8_1  (
            .in0(N__16937),
            .in1(N__17039),
            .in2(N__16998),
            .in3(N__19588),
            .lcout(\Lab_UT.N_65 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Mtens_alarm.q_RNI7VK11_3_LC_7_8_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mtens_alarm.q_RNI7VK11_3_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Mtens_alarm.q_RNI7VK11_3_LC_7_8_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Lab_UT.didp.Mtens_alarm.q_RNI7VK11_3_LC_7_8_2  (
            .in0(N__26833),
            .in1(N__25533),
            .in2(_gnd_net_),
            .in3(N__19664),
            .lcout(\Lab_UT.Mten_at_3 ),
            .ltout(\Lab_UT.Mten_at_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment4.segment_1_3_LC_7_8_3 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment4.segment_1_3_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment4.segment_1_3_LC_7_8_3 .LUT_INIT=16'b1101110011011111;
    LogicCell40 \Lab_UT.bcd2segment4.segment_1_3_LC_7_8_3  (
            .in0(N__16858),
            .in1(N__17038),
            .in2(N__16873),
            .in3(N__16833),
            .lcout(\Lab_UT.segment_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment4.segmentUQ_0_o2_5_LC_7_8_4 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment4.segmentUQ_0_o2_5_LC_7_8_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment4.segmentUQ_0_o2_5_LC_7_8_4 .LUT_INIT=16'b0001110100000000;
    LogicCell40 \Lab_UT.bcd2segment4.segmentUQ_0_o2_5_LC_7_8_4  (
            .in0(N__25852),
            .in1(N__19665),
            .in2(N__26890),
            .in3(N__16935),
            .lcout(\Lab_UT.N_69_0 ),
            .ltout(\Lab_UT.N_69_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment4.segmentUQ_i_a3_0_2_LC_7_8_5 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment4.segmentUQ_i_a3_0_2_LC_7_8_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment4.segmentUQ_i_a3_0_2_LC_7_8_5 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \Lab_UT.bcd2segment4.segmentUQ_i_a3_0_2_LC_7_8_5  (
            .in0(N__16983),
            .in1(_gnd_net_),
            .in2(N__16849),
            .in3(N__17037),
            .lcout(\Lab_UT.N_92 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment4.segmentUQ_0_o3_5_LC_7_8_6 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment4.segmentUQ_0_o3_5_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment4.segmentUQ_0_o3_5_LC_7_8_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Lab_UT.bcd2segment4.segmentUQ_0_o3_5_LC_7_8_6  (
            .in0(_gnd_net_),
            .in1(N__19587),
            .in2(_gnd_net_),
            .in3(N__16934),
            .lcout(\Lab_UT.N_67_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment4.segmentUQ_i_a3_2_LC_7_8_7 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment4.segmentUQ_i_a3_2_LC_7_8_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment4.segmentUQ_i_a3_2_LC_7_8_7 .LUT_INIT=16'b1011000000000000;
    LogicCell40 \Lab_UT.bcd2segment4.segmentUQ_i_a3_2_LC_7_8_7  (
            .in0(N__16936),
            .in1(N__17033),
            .in2(N__16999),
            .in3(N__19589),
            .lcout(\Lab_UT.N_91 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment4.segmentUQ_i_a4_3_LC_7_9_0 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment4.segmentUQ_i_a4_3_LC_7_9_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment4.segmentUQ_i_a4_3_LC_7_9_0 .LUT_INIT=16'b1000100000100010;
    LogicCell40 \Lab_UT.bcd2segment4.segmentUQ_i_a4_3_LC_7_9_0  (
            .in0(N__17032),
            .in1(N__19590),
            .in2(_gnd_net_),
            .in3(N__16938),
            .lcout(\Lab_UT.N_83 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Mtens_alarm.q_RNI1PK11_0_LC_7_9_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mtens_alarm.q_RNI1PK11_0_LC_7_9_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Mtens_alarm.q_RNI1PK11_0_LC_7_9_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Lab_UT.didp.Mtens_alarm.q_RNI1PK11_0_LC_7_9_1  (
            .in0(N__30038),
            .in1(N__25061),
            .in2(_gnd_net_),
            .in3(N__19645),
            .lcout(\Lab_UT.Mten_at_0 ),
            .ltout(\Lab_UT.Mten_at_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment4.segmentUQ_i_a3_0_4_LC_7_9_2 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment4.segmentUQ_i_a3_0_4_LC_7_9_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment4.segmentUQ_i_a3_0_4_LC_7_9_2 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \Lab_UT.bcd2segment4.segmentUQ_i_a3_0_4_LC_7_9_2  (
            .in0(N__16987),
            .in1(_gnd_net_),
            .in2(N__16951),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.N_77 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Mtens_alarm.q_RNI3RK11_1_LC_7_9_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mtens_alarm.q_RNI3RK11_1_LC_7_9_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Mtens_alarm.q_RNI3RK11_1_LC_7_9_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Lab_UT.didp.Mtens_alarm.q_RNI3RK11_1_LC_7_9_3  (
            .in0(N__27948),
            .in1(N__26354),
            .in2(_gnd_net_),
            .in3(N__19644),
            .lcout(\Lab_UT.Mten_at_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Mtens_alarm.q_0_LC_7_9_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mtens_alarm.q_0_LC_7_9_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.Mtens_alarm.q_0_LC_7_9_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \Lab_UT.didp.Mtens_alarm.q_0_LC_7_9_4  (
            .in0(N__25062),
            .in1(N__23014),
            .in2(_gnd_net_),
            .in3(N__29102),
            .lcout(\Lab_UT.di_AMtens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29401),
            .ce(),
            .sr(N__26065));
    defparam \Lab_UT.didp.Mtens_alarm.q_1_LC_7_9_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mtens_alarm.q_1_LC_7_9_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.Mtens_alarm.q_1_LC_7_9_5 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \Lab_UT.didp.Mtens_alarm.q_1_LC_7_9_5  (
            .in0(N__28821),
            .in1(_gnd_net_),
            .in2(N__23020),
            .in3(N__26355),
            .lcout(\Lab_UT.di_AMtens_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29401),
            .ce(),
            .sr(N__26065));
    defparam \Lab_UT.dictrl.currState_2_2_LC_7_9_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_2_LC_7_9_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.currState_2_2_LC_7_9_6 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \Lab_UT.dictrl.currState_2_2_LC_7_9_6  (
            .in0(N__17725),
            .in1(N__17419),
            .in2(N__17083),
            .in3(N__17401),
            .lcout(\Lab_UT.dictrl.currStateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29401),
            .ce(),
            .sr(N__26065));
    defparam \Lab_UT.dictrl.currState_0_ret_14_LC_7_10_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_14_LC_7_10_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.currState_0_ret_14_LC_7_10_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_14_LC_7_10_0  (
            .in0(N__21520),
            .in1(N__20653),
            .in2(N__20815),
            .in3(N__21034),
            .lcout(\Lab_UT.dictrl.un2_dicAlarmTrig ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29395),
            .ce(),
            .sr(N__26067));
    defparam \Lab_UT.dictrl.currState_0_ret_3_LC_7_10_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_3_LC_7_10_1 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.currState_0_ret_3_LC_7_10_1 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_3_LC_7_10_1  (
            .in0(N__21033),
            .in1(N__21521),
            .in2(N__20794),
            .in3(N__20634),
            .lcout(\Lab_UT.dictrl.r_Sone_init5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29395),
            .ce(),
            .sr(N__26067));
    defparam \Lab_UT.dictrl.currState_0_ret_29_RNO_0_LC_7_10_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_29_RNO_0_LC_7_10_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_0_ret_29_RNO_0_LC_7_10_2 .LUT_INIT=16'b0110101011101011;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_29_RNO_0_LC_7_10_2  (
            .in0(N__21519),
            .in1(N__21032),
            .in2(N__20659),
            .in3(N__20747),
            .lcout(\Lab_UT.dictrl.g0_13_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_RNII4T093_0_2_LC_7_10_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_RNII4T093_0_2_LC_7_10_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_RNII4T093_0_2_LC_7_10_3 .LUT_INIT=16'b0110110011001101;
    LogicCell40 \Lab_UT.dictrl.currState_2_RNII4T093_0_2_LC_7_10_3  (
            .in0(N__21028),
            .in1(N__21515),
            .in2(N__20792),
            .in3(N__20623),
            .lcout(\Lab_UT.dictrl.g0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_RNO_10_1_LC_7_10_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_RNO_10_1_LC_7_10_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_RNO_10_1_LC_7_10_4 .LUT_INIT=16'b0100101000001010;
    LogicCell40 \Lab_UT.dictrl.nextState_RNO_10_1_LC_7_10_4  (
            .in0(N__21516),
            .in1(N__21030),
            .in2(N__20657),
            .in3(N__20742),
            .lcout(\Lab_UT.dictrl.g0_i_o4_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_RNII4T093_1_2_LC_7_10_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_RNII4T093_1_2_LC_7_10_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_RNII4T093_1_2_LC_7_10_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \Lab_UT.dictrl.currState_2_RNII4T093_1_2_LC_7_10_5  (
            .in0(N__21029),
            .in1(N__21517),
            .in2(N__20793),
            .in3(N__20627),
            .lcout(\Lab_UT.dictrl.r_dicLdMtens16_reti ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_RNII4T093_2_LC_7_10_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_RNII4T093_2_LC_7_10_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_RNII4T093_2_LC_7_10_6 .LUT_INIT=16'b0110101110101011;
    LogicCell40 \Lab_UT.dictrl.currState_2_RNII4T093_2_LC_7_10_6  (
            .in0(N__21518),
            .in1(N__21031),
            .in2(N__20658),
            .in3(N__20746),
            .lcout(\Lab_UT.dictrl.currState_0_ret_20and_1_0 ),
            .ltout(\Lab_UT.dictrl.currState_0_ret_20and_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_RNI82L3I6_2_LC_7_10_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_RNI82L3I6_2_LC_7_10_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_RNI82L3I6_2_LC_7_10_7 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \Lab_UT.dictrl.currState_2_RNI82L3I6_2_LC_7_10_7  (
            .in0(N__24689),
            .in1(_gnd_net_),
            .in2(N__17116),
            .in3(N__20118),
            .lcout(\Lab_UT.dictrl.N_258_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.dicLdASones_RNI1C3E5_LC_7_11_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.dicLdASones_RNI1C3E5_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.dicLdASones_RNI1C3E5_LC_7_11_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \Lab_UT.dictrl.dicLdASones_RNI1C3E5_LC_7_11_0  (
            .in0(N__17364),
            .in1(N__20506),
            .in2(_gnd_net_),
            .in3(N__17374),
            .lcout(\Lab_UT.ld_enable_ASones ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_3_3_rep1_RNI2J197_LC_7_11_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_3_3_rep1_RNI2J197_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_3_3_rep1_RNI2J197_LC_7_11_2 .LUT_INIT=16'b1010110010100000;
    LogicCell40 \Lab_UT.dictrl.currState_3_3_rep1_RNI2J197_LC_7_11_2  (
            .in0(N__17113),
            .in1(N__27802),
            .in2(N__20396),
            .in3(N__27544),
            .lcout(\Lab_UT.dictrl.N_13 ),
            .ltout(\Lab_UT.dictrl.N_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_3_3_rep1_RNIKKEKM_LC_7_11_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_3_3_rep1_RNIKKEKM_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_3_3_rep1_RNIKKEKM_LC_7_11_3 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \Lab_UT.dictrl.currState_3_3_rep1_RNIKKEKM_LC_7_11_3  (
            .in0(N__17724),
            .in1(N__17415),
            .in2(N__17404),
            .in3(N__17394),
            .lcout(\Lab_UT.dictrl.nextStateZ0Z_2 ),
            .ltout(\Lab_UT.dictrl.nextStateZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_3_3_rep1_RNI39J171_LC_7_11_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_3_3_rep1_RNI39J171_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_3_3_rep1_RNI39J171_LC_7_11_4 .LUT_INIT=16'b0000000000001010;
    LogicCell40 \Lab_UT.dictrl.currState_3_3_rep1_RNI39J171_LC_7_11_4  (
            .in0(N__21514),
            .in1(_gnd_net_),
            .in2(N__17377),
            .in3(N__24679),
            .lcout(\Lab_UT.dictrl.currState_ret_1and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_RNIMNQP4_2_LC_7_11_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_RNIMNQP4_2_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_RNIMNQP4_2_LC_7_11_5 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \Lab_UT.dictrl.currState_2_RNIMNQP4_2_LC_7_11_5  (
            .in0(N__27545),
            .in1(_gnd_net_),
            .in2(N__27814),
            .in3(N__23670),
            .lcout(\Lab_UT.dictrl.dicLdASones_rst ),
            .ltout(\Lab_UT.dictrl.dicLdASones_rst_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.dicLdASones_LC_7_11_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.dicLdASones_LC_7_11_6 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.dictrl.dicLdASones_LC_7_11_6 .LUT_INIT=16'b1010101011100010;
    LogicCell40 \Lab_UT.dictrl.dicLdASones_LC_7_11_6  (
            .in0(N__17365),
            .in1(N__20507),
            .in2(N__17368),
            .in3(N__20560),
            .lcout(\Lab_UT.dictrl.dicLdASonesZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29391),
            .ce(),
            .sr(N__23671));
    defparam \Lab_UT.dictrl.currState_2_RNIFK4DG_1_LC_7_11_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_RNIFK4DG_1_LC_7_11_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_RNIFK4DG_1_LC_7_11_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.dictrl.currState_2_RNIFK4DG_1_LC_7_11_7  (
            .in0(_gnd_net_),
            .in1(N__24676),
            .in2(_gnd_net_),
            .in3(N__21513),
            .lcout(\Lab_UT.dictrl.N_5ctr ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_0_ret_1_LC_7_12_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_1_LC_7_12_0 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.currState_0_ret_1_LC_7_12_0 .LUT_INIT=16'b1010001000000010;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_1_LC_7_12_0  (
            .in0(N__21040),
            .in1(N__17308),
            .in2(N__17185),
            .in3(N__17266),
            .lcout(\Lab_UT.dictrl.r_Sone_init5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29385),
            .ce(),
            .sr(N__26070));
    defparam \Lab_UT.dictrl.currState_0_ret_5_LC_7_12_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_5_LC_7_12_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.currState_0_ret_5_LC_7_12_1 .LUT_INIT=16'b0000000000111010;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_5_LC_7_12_1  (
            .in0(N__17307),
            .in1(N__17265),
            .in2(N__17183),
            .in3(N__21041),
            .lcout(\Lab_UT.dictrl.r_dicLdMtens14_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29385),
            .ce(),
            .sr(N__26070));
    defparam \Lab_UT.dictrl.currState_2_RNIRPGDN_1_LC_7_12_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_RNIRPGDN_1_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_RNIRPGDN_1_LC_7_12_2 .LUT_INIT=16'b1110110011101111;
    LogicCell40 \Lab_UT.dictrl.currState_2_RNIRPGDN_1_LC_7_12_2  (
            .in0(N__17264),
            .in1(N__24684),
            .in2(N__17184),
            .in3(N__17306),
            .lcout(\Lab_UT.dictrl.N_7ctr ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_RNI4F3LS1_1_LC_7_12_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_RNI4F3LS1_1_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_RNI4F3LS1_1_LC_7_12_3 .LUT_INIT=16'b0011101000000000;
    LogicCell40 \Lab_UT.dictrl.currState_2_RNI4F3LS1_1_LC_7_12_3  (
            .in0(N__17305),
            .in1(N__17263),
            .in2(N__17182),
            .in3(N__21038),
            .lcout(\Lab_UT.dictrl.r_dicLdMtens15_1i ),
            .ltout(\Lab_UT.dictrl.r_dicLdMtens15_1i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_RNI7OMM33_1_LC_7_12_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_RNI7OMM33_1_LC_7_12_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_RNI7OMM33_1_LC_7_12_4 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Lab_UT.dictrl.currState_2_RNI7OMM33_1_LC_7_12_4  (
            .in0(N__21574),
            .in1(N__24685),
            .in2(N__17602),
            .in3(N__20757),
            .lcout(\Lab_UT.dictrl.currState_ret_3and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_0_ret_28_RNO_3_LC_7_12_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_28_RNO_3_LC_7_12_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_0_ret_28_RNO_3_LC_7_12_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_28_RNO_3_LC_7_12_5  (
            .in0(N__20756),
            .in1(N__21573),
            .in2(_gnd_net_),
            .in3(N__21039),
            .lcout(),
            .ltout(\Lab_UT.dictrl.currState_0_ret_28_RNOZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_0_ret_28_RNO_1_LC_7_12_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_28_RNO_1_LC_7_12_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_0_ret_28_RNO_1_LC_7_12_6 .LUT_INIT=16'b0010011110101111;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_28_RNO_1_LC_7_12_6  (
            .in0(N__17587),
            .in1(N__17571),
            .in2(N__17491),
            .in3(N__17479),
            .lcout(\Lab_UT.dictrl.N_8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_RNIS2IML1_2_LC_7_12_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_RNIS2IML1_2_LC_7_12_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_RNIS2IML1_2_LC_7_12_7 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \Lab_UT.dictrl.currState_2_RNIS2IML1_2_LC_7_12_7  (
            .in0(N__24683),
            .in1(N__21572),
            .in2(_gnd_net_),
            .in3(N__21037),
            .lcout(\Lab_UT.dictrl.r_dicLdMtens21_1_reti ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.decoder.g0_10_LC_7_13_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.decoder.g0_10_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.decoder.g0_10_LC_7_13_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.decoder.g0_10_LC_7_13_0  (
            .in0(N__17710),
            .in1(N__17472),
            .in2(N__18186),
            .in3(N__17660),
            .lcout(),
            .ltout(\Lab_UT.dictrl.de_littleA_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_3_LC_7_13_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_3_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_3_LC_7_13_1 .LUT_INIT=16'b0000001000001010;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__g0_3_LC_7_13_1  (
            .in0(N__20891),
            .in1(N__24217),
            .in2(N__17458),
            .in3(N__27748),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_37_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_RNIQ4BA8_1_LC_7_13_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_RNIQ4BA8_1_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_RNIQ4BA8_1_LC_7_13_2 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \Lab_UT.dictrl.currState_2_RNIQ4BA8_1_LC_7_13_2  (
            .in0(N__17926),
            .in1(N__18070),
            .in2(N__17455),
            .in3(N__18055),
            .lcout(\Lab_UT.dictrl.g0_15_rn_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_3_3_rep1_RNIRM2Q_LC_7_13_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_3_3_rep1_RNIRM2Q_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_3_3_rep1_RNIRM2Q_LC_7_13_3 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \Lab_UT.dictrl.currState_3_3_rep1_RNIRM2Q_LC_7_13_3  (
            .in0(N__20394),
            .in1(N__25025),
            .in2(N__23458),
            .in3(N__17925),
            .lcout(\Lab_UT.dictrl.G_19_0_a7_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_2_rep1_es_RNIELCR_LC_7_13_4 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_2_rep1_es_RNIELCR_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_2_rep1_es_RNIELCR_LC_7_13_4 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \buart.Z_rx.bitcount_2_rep1_es_RNIELCR_LC_7_13_4  (
            .in0(N__21703),
            .in1(N__21937),
            .in2(N__21780),
            .in3(N__17697),
            .lcout(G_19_0_a7_4_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_RNIEPCJ_1_LC_7_13_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_RNIEPCJ_1_LC_7_13_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_RNIEPCJ_1_LC_7_13_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.dictrl.currState_2_RNIEPCJ_1_LC_7_13_5  (
            .in0(_gnd_net_),
            .in1(N__18053),
            .in2(_gnd_net_),
            .in3(N__17924),
            .lcout(\Lab_UT.dictrl.currState_2_RNIEPCJZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_RNI2SKC_3_LC_7_13_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_RNI2SKC_3_LC_7_13_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_RNI2SKC_3_LC_7_13_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Lab_UT.dictrl.nextState_RNI2SKC_3_LC_7_13_6  (
            .in0(N__18088),
            .in1(N__23448),
            .in2(_gnd_net_),
            .in3(N__20393),
            .lcout(\Lab_UT.dictrl.N_1612_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_RNIEGFT_0_LC_7_13_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_RNIEGFT_0_LC_7_13_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_RNIEGFT_0_LC_7_13_7 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Lab_UT.dictrl.currState_2_RNIEGFT_0_LC_7_13_7  (
            .in0(N__23452),
            .in1(N__18054),
            .in2(N__21268),
            .in3(N__17927),
            .lcout(\Lab_UT.dictrl.G_19_0_a7_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.decoder.g0_2_2_LC_7_14_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.decoder.g0_2_2_LC_7_14_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.decoder.g0_2_2_LC_7_14_0 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \Lab_UT.dictrl.decoder.g0_2_2_LC_7_14_0  (
            .in0(N__21832),
            .in1(N__21918),
            .in2(N__21991),
            .in3(N__17695),
            .lcout(\Lab_UT.dictrl.decoder.g0_2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.decoder.de_cr_2_LC_7_14_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.decoder.de_cr_2_LC_7_14_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.decoder.de_cr_2_LC_7_14_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.dictrl.decoder.de_cr_2_LC_7_14_1  (
            .in0(_gnd_net_),
            .in1(N__21891),
            .in2(_gnd_net_),
            .in3(N__17616),
            .lcout(Lab_UT_dictrl_decoder_de_cr_2),
            .ltout(Lab_UT_dictrl_decoder_de_cr_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.decoder.g0_4_3_LC_7_14_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.decoder.g0_4_3_LC_7_14_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.decoder.g0_4_3_LC_7_14_2 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \Lab_UT.dictrl.decoder.g0_4_3_LC_7_14_2  (
            .in0(N__21833),
            .in1(_gnd_net_),
            .in2(N__17701),
            .in3(N__17696),
            .lcout(),
            .ltout(\Lab_UT.dictrl.decoder.g0_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.decoder.g0_11_LC_7_14_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.decoder.g0_11_LC_7_14_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.decoder.g0_11_LC_7_14_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.decoder.g0_11_LC_7_14_3  (
            .in0(N__21358),
            .in1(N__18172),
            .in2(N__17671),
            .in3(N__17667),
            .lcout(\Lab_UT.dictrl.de_cr_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_fast_2_LC_7_14_4 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_2_LC_7_14_4 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_fast_2_LC_7_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_fast_2_LC_7_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28906),
            .lcout(bu_rx_data_fast_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29377),
            .ce(N__25423),
            .sr(N__26097));
    defparam \buart.Z_rx.shifter_fast_1_LC_7_14_7 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_1_LC_7_14_7 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_fast_1_LC_7_14_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_fast_1_LC_7_14_7  (
            .in0(N__28573),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_fast_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29377),
            .ce(N__25423),
            .sr(N__26097));
    defparam \Lab_UT.dictrl.decoder.g0_13_LC_7_15_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.decoder.g0_13_LC_7_15_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.decoder.g0_13_LC_7_15_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.decoder.g0_13_LC_7_15_0  (
            .in0(N__18175),
            .in1(N__18409),
            .in2(N__18331),
            .in3(N__18367),
            .lcout(\Lab_UT.dictrl.de_cr_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.decoder.de_cr_1_1_LC_7_15_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.decoder.de_cr_1_1_LC_7_15_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.decoder.de_cr_1_1_LC_7_15_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Lab_UT.dictrl.decoder.de_cr_1_1_LC_7_15_1  (
            .in0(N__24441),
            .in1(N__25300),
            .in2(N__24294),
            .in3(N__21414),
            .lcout(Lab_UT_dictrl_decoder_de_cr_1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.decoder.g0_17_LC_7_15_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.decoder.g0_17_LC_7_15_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.decoder.g0_17_LC_7_15_2 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \Lab_UT.dictrl.decoder.g0_17_LC_7_15_2  (
            .in0(N__25374),
            .in1(N__18307),
            .in2(N__29048),
            .in3(N__18273),
            .lcout(\Lab_UT.dictrl.decoder.g0_4Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.decoder.g0_16_LC_7_15_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.decoder.g0_16_LC_7_15_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.decoder.g0_16_LC_7_15_3 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \Lab_UT.dictrl.decoder.g0_16_LC_7_15_3  (
            .in0(N__28597),
            .in1(N__28924),
            .in2(_gnd_net_),
            .in3(N__18226),
            .lcout(),
            .ltout(\Lab_UT.dictrl.decoder.g0_3_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.decoder.g0_15_LC_7_15_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.decoder.g0_15_LC_7_15_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.decoder.g0_15_LC_7_15_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.decoder.g0_15_LC_7_15_4  (
            .in0(N__18174),
            .in1(N__18385),
            .in2(N__18379),
            .in3(N__18366),
            .lcout(\Lab_UT.dictrl.de_cr_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.decoder.g0_14_LC_7_15_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.decoder.g0_14_LC_7_15_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.decoder.g0_14_LC_7_15_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Lab_UT.dictrl.decoder.g0_14_LC_7_15_5  (
            .in0(N__18274),
            .in1(N__25375),
            .in2(N__18320),
            .in3(N__29026),
            .lcout(\Lab_UT.dictrl.decoder.g0_4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_15_LC_7_15_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_15_LC_7_15_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_15_LC_7_15_6 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__g0_15_LC_7_15_6  (
            .in0(N__25373),
            .in1(N__18306),
            .in2(N__29047),
            .in3(N__18272),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_12_LC_7_15_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_12_LC_7_15_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_12_LC_7_15_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__g0_12_LC_7_15_7  (
            .in0(N__24442),
            .in1(N__18225),
            .in2(N__18190),
            .in3(N__18173),
            .lcout(\Lab_UT.dictrl.g0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.uu0.l_count_6_LC_8_1_0 .C_ON=1'b0;
    defparam \Lab_UT.uu0.l_count_6_LC_8_1_0 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.uu0.l_count_6_LC_8_1_0 .LUT_INIT=16'b0001010101000000;
    LogicCell40 \Lab_UT.uu0.l_count_6_LC_8_1_0  (
            .in0(N__23233),
            .in1(N__22194),
            .in2(N__18517),
            .in3(N__22036),
            .lcout(\Lab_UT.uu0.l_countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29471),
            .ce(N__22173),
            .sr(N__26102));
    defparam \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_8_1_1 .C_ON=1'b0;
    defparam \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_8_1_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_8_1_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_8_1_1  (
            .in0(N__22035),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18513),
            .lcout(),
            .ltout(\Lab_UT.uu0.un99_ci_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.uu0.l_count_7_LC_8_1_2 .C_ON=1'b0;
    defparam \Lab_UT.uu0.l_count_7_LC_8_1_2 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.uu0.l_count_7_LC_8_1_2 .LUT_INIT=16'b0001010101000000;
    LogicCell40 \Lab_UT.uu0.l_count_7_LC_8_1_2  (
            .in0(N__23234),
            .in1(N__22195),
            .in2(N__18520),
            .in3(N__18502),
            .lcout(\Lab_UT.uu0.l_countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29471),
            .ce(N__22173),
            .sr(N__26102));
    defparam \Lab_UT.uu0.l_count_16_LC_8_1_3 .C_ON=1'b0;
    defparam \Lab_UT.uu0.l_count_16_LC_8_1_3 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.uu0.l_count_16_LC_8_1_3 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \Lab_UT.uu0.l_count_16_LC_8_1_3  (
            .in0(N__18621),
            .in1(N__22578),
            .in2(N__18609),
            .in3(N__23232),
            .lcout(\Lab_UT.uu0.l_countZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29471),
            .ce(N__22173),
            .sr(N__26102));
    defparam \Lab_UT.uu0.l_count_17_LC_8_1_4 .C_ON=1'b0;
    defparam \Lab_UT.uu0.l_count_17_LC_8_1_4 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.uu0.l_count_17_LC_8_1_4 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \Lab_UT.uu0.l_count_17_LC_8_1_4  (
            .in0(N__22579),
            .in1(N__18601),
            .in2(N__18486),
            .in3(N__18622),
            .lcout(\Lab_UT.uu0.l_countZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29471),
            .ce(N__22173),
            .sr(N__26102));
    defparam \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_8_1_5 .C_ON=1'b0;
    defparam \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_8_1_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_8_1_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_8_1_5  (
            .in0(_gnd_net_),
            .in1(N__22214),
            .in2(_gnd_net_),
            .in3(N__22128),
            .lcout(\Lab_UT.uu0.un88_ci_3 ),
            .ltout(\Lab_UT.uu0.un88_ci_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_8_1_6 .C_ON=1'b0;
    defparam \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_8_1_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_8_1_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_8_1_6  (
            .in0(N__22192),
            .in1(N__22034),
            .in2(N__18505),
            .in3(N__18501),
            .lcout(\Lab_UT.uu0.un110_ci ),
            .ltout(\Lab_UT.uu0.un110_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_8_1_7 .C_ON=1'b0;
    defparam \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_8_1_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_8_1_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_8_1_7  (
            .in0(N__18620),
            .in1(N__18479),
            .in2(N__18463),
            .in3(N__22577),
            .lcout(\Lab_UT.uu0.un220_ci ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.uu0.l_count_10_LC_8_2_0 .C_ON=1'b0;
    defparam \Lab_UT.uu0.l_count_10_LC_8_2_0 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.uu0.l_count_10_LC_8_2_0 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \Lab_UT.uu0.l_count_10_LC_8_2_0  (
            .in0(N__18555),
            .in1(N__18454),
            .in2(N__18608),
            .in3(N__18428),
            .lcout(\Lab_UT.uu0.l_countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29464),
            .ce(N__22170),
            .sr(N__26100));
    defparam \Lab_UT.uu0.l_count_RNIKE6P_2_LC_8_2_1 .C_ON=1'b0;
    defparam \Lab_UT.uu0.l_count_RNIKE6P_2_LC_8_2_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.uu0.l_count_RNIKE6P_2_LC_8_2_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Lab_UT.uu0.l_count_RNIKE6P_2_LC_8_2_1  (
            .in0(N__18427),
            .in1(N__18554),
            .in2(N__18671),
            .in3(N__22235),
            .lcout(),
            .ltout(\Lab_UT.uu0.un4_l_count_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.uu0.l_count_RNIAK6Q1_4_LC_8_2_2 .C_ON=1'b0;
    defparam \Lab_UT.uu0.l_count_RNIAK6Q1_4_LC_8_2_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.uu0.l_count_RNIAK6Q1_4_LC_8_2_2 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \Lab_UT.uu0.l_count_RNIAK6Q1_4_LC_8_2_2  (
            .in0(N__25200),
            .in1(N__22213),
            .in2(N__18700),
            .in3(N__18643),
            .lcout(\Lab_UT.uu0.un4_l_count_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.uu0.l_count_14_LC_8_2_3 .C_ON=1'b0;
    defparam \Lab_UT.uu0.l_count_14_LC_8_2_3 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.uu0.l_count_14_LC_8_2_3 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \Lab_UT.uu0.l_count_14_LC_8_2_3  (
            .in0(N__18690),
            .in1(N__18646),
            .in2(N__18672),
            .in3(N__18593),
            .lcout(\Lab_UT.uu0.l_countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29464),
            .ce(N__22170),
            .sr(N__26100));
    defparam \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_8_2_4 .C_ON=1'b0;
    defparam \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_8_2_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_8_2_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_8_2_4  (
            .in0(N__18670),
            .in1(N__18689),
            .in2(_gnd_net_),
            .in3(N__18645),
            .lcout(),
            .ltout(\Lab_UT.uu0.un187_ci_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.uu0.l_count_15_LC_8_2_5 .C_ON=1'b0;
    defparam \Lab_UT.uu0.l_count_15_LC_8_2_5 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.uu0.l_count_15_LC_8_2_5 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \Lab_UT.uu0.l_count_15_LC_8_2_5  (
            .in0(N__22057),
            .in1(N__18594),
            .in2(N__18697),
            .in3(N__23223),
            .lcout(\Lab_UT.uu0.l_countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29464),
            .ce(N__22170),
            .sr(N__26100));
    defparam \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_8_2_6 .C_ON=1'b0;
    defparam \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_8_2_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_8_2_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_8_2_6  (
            .in0(N__22056),
            .in1(N__18688),
            .in2(N__18673),
            .in3(N__18644),
            .lcout(\Lab_UT.uu0.un198_ci_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.uu0.l_count_8_LC_8_2_7 .C_ON=1'b0;
    defparam \Lab_UT.uu0.l_count_8_LC_8_2_7 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.uu0.l_count_8_LC_8_2_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Lab_UT.uu0.l_count_8_LC_8_2_7  (
            .in0(_gnd_net_),
            .in1(N__18592),
            .in2(_gnd_net_),
            .in3(N__18556),
            .lcout(\Lab_UT.uu0.l_countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29464),
            .ce(N__22170),
            .sr(N__26100));
    defparam \uu2.w_addr_user_RNI0FES5_2_LC_8_3_0 .C_ON=1'b0;
    defparam \uu2.w_addr_user_RNI0FES5_2_LC_8_3_0 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_RNI0FES5_2_LC_8_3_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \uu2.w_addr_user_RNI0FES5_2_LC_8_3_0  (
            .in0(_gnd_net_),
            .in1(N__22312),
            .in2(_gnd_net_),
            .in3(N__22423),
            .lcout(\uu2.un28_w_addr_user_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un1_w_user_lf_LC_8_3_1 .C_ON=1'b0;
    defparam \uu2.un1_w_user_lf_LC_8_3_1 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_w_user_lf_LC_8_3_1 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \uu2.un1_w_user_lf_LC_8_3_1  (
            .in0(N__18823),
            .in1(N__22280),
            .in2(N__25687),
            .in3(N__22827),
            .lcout(\uu2.un1_w_user_lf_0 ),
            .ltout(\uu2.un1_w_user_lf_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_RNIMJ3O2_2_LC_8_3_2 .C_ON=1'b0;
    defparam \uu2.w_addr_user_RNIMJ3O2_2_LC_8_3_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_RNIMJ3O2_2_LC_8_3_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \uu2.w_addr_user_RNIMJ3O2_2_LC_8_3_2  (
            .in0(N__18891),
            .in1(N__26143),
            .in2(N__18523),
            .in3(N__18879),
            .lcout(\uu2.w_addr_user_RNIMJ3O2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vram_wr_en_0_i_LC_8_3_3 .C_ON=1'b0;
    defparam \uu2.vram_wr_en_0_i_LC_8_3_3 .SEQ_MODE=4'b0000;
    defparam \uu2.vram_wr_en_0_i_LC_8_3_3 .LUT_INIT=16'b0111011100110011;
    LogicCell40 \uu2.vram_wr_en_0_i_LC_8_3_3  (
            .in0(N__18880),
            .in1(N__29490),
            .in2(_gnd_net_),
            .in3(N__22294),
            .lcout(\uu2.vram_wr_en_0_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_RNIARA43_2_LC_8_3_4 .C_ON=1'b0;
    defparam \uu2.w_addr_user_RNIARA43_2_LC_8_3_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_RNIARA43_2_LC_8_3_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \uu2.w_addr_user_RNIARA43_2_LC_8_3_4  (
            .in0(N__22293),
            .in1(N__18898),
            .in2(N__18892),
            .in3(N__18878),
            .lcout(\uu2.un28_w_addr_user_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un1_w_user_cr_LC_8_3_5 .C_ON=1'b0;
    defparam \uu2.un1_w_user_cr_LC_8_3_5 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_w_user_cr_LC_8_3_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \uu2.un1_w_user_cr_LC_8_3_5  (
            .in0(N__25683),
            .in1(N__18829),
            .in2(N__25594),
            .in3(N__22661),
            .lcout(\uu2.un1_w_user_cr_0 ),
            .ltout(\uu2.un1_w_user_cr_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un4_w_user_data_rdy_0_LC_8_3_6 .C_ON=1'b0;
    defparam \uu2.un4_w_user_data_rdy_0_LC_8_3_6 .SEQ_MODE=4'b0000;
    defparam \uu2.un4_w_user_data_rdy_0_LC_8_3_6 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \uu2.un4_w_user_data_rdy_0_LC_8_3_6  (
            .in0(N__22292),
            .in1(_gnd_net_),
            .in2(N__18868),
            .in3(_gnd_net_),
            .lcout(\uu2.un4_w_user_data_rdyZ0Z_0 ),
            .ltout(\uu2.un4_w_user_data_rdyZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_14_LC_8_3_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_14_LC_8_3_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_14_LC_8_3_7 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_14_LC_8_3_7  (
            .in0(_gnd_net_),
            .in1(N__18863),
            .in2(N__18847),
            .in3(N__22281),
            .lcout(\uu2.mem0.w_data_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un1_w_user_cr_4_LC_8_4_0 .C_ON=1'b0;
    defparam \uu2.un1_w_user_cr_4_LC_8_4_0 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_w_user_cr_4_LC_8_4_0 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \uu2.un1_w_user_cr_4_LC_8_4_0  (
            .in0(N__22613),
            .in1(N__22632),
            .in2(N__22282),
            .in3(N__22820),
            .lcout(\uu2.un1_w_user_crZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un1_w_user_lf_4_LC_8_4_1 .C_ON=1'b0;
    defparam \uu2.un1_w_user_lf_4_LC_8_4_1 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_w_user_lf_4_LC_8_4_1 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \uu2.un1_w_user_lf_4_LC_8_4_1  (
            .in0(N__22631),
            .in1(N__25586),
            .in2(N__22665),
            .in3(N__22614),
            .lcout(\uu2.un1_w_user_lfZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_10_LC_8_4_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_10_LC_8_4_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_10_LC_8_4_2 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_10_LC_8_4_2  (
            .in0(N__18751),
            .in1(N__25590),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uu2.mem0.w_data_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_LC_8_4_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_LC_8_4_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_LC_8_4_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_LC_8_4_3  (
            .in0(N__19062),
            .in1(N__18750),
            .in2(_gnd_net_),
            .in3(N__19495),
            .lcout(\uu2.mem0.w_addr_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_0_LC_8_4_4 .C_ON=1'b0;
    defparam \uu2.w_addr_user_0_LC_8_4_4 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_0_LC_8_4_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.w_addr_user_0_LC_8_4_4  (
            .in0(_gnd_net_),
            .in1(N__19064),
            .in2(_gnd_net_),
            .in3(N__22424),
            .lcout(\uu2.w_addr_userZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_0C_net ),
            .ce(),
            .sr(N__22327));
    defparam \uu2.w_addr_user_1_LC_8_4_5 .C_ON=1'b0;
    defparam \uu2.w_addr_user_1_LC_8_4_5 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_1_LC_8_4_5 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \uu2.w_addr_user_1_LC_8_4_5  (
            .in0(N__22425),
            .in1(_gnd_net_),
            .in2(N__19069),
            .in3(N__18968),
            .lcout(\uu2.w_addr_userZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_0C_net ),
            .ce(),
            .sr(N__22327));
    defparam \uu2.w_addr_user_2_LC_8_4_6 .C_ON=1'b0;
    defparam \uu2.w_addr_user_2_LC_8_4_6 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_2_LC_8_4_6 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.w_addr_user_2_LC_8_4_6  (
            .in0(N__18969),
            .in1(N__19068),
            .in2(N__19034),
            .in3(N__22426),
            .lcout(\uu2.w_addr_userZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_0C_net ),
            .ce(),
            .sr(N__22327));
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_4__un404_ci_LC_8_4_7 .C_ON=1'b0;
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_4__un404_ci_LC_8_4_7 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_4__un404_ci_LC_8_4_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.vbuf_w_addr_user.counter_gen_label_4__un404_ci_LC_8_4_7  (
            .in0(N__19063),
            .in1(N__19023),
            .in2(N__18997),
            .in3(N__18967),
            .lcout(\uu2.un404_ci ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.curr_LED_1_LC_8_5_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.curr_LED_1_LC_8_5_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.curr_LED_1_LC_8_5_0 .LUT_INIT=16'b0001010101000000;
    LogicCell40 \Lab_UT.didp.curr_LED_1_LC_8_5_0  (
            .in0(N__26151),
            .in1(N__29725),
            .in2(N__25456),
            .in3(N__29612),
            .lcout(\Lab_UT.didp.curr_LEDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29441),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.curr_LED_0_LC_8_5_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.curr_LED_0_LC_8_5_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.curr_LED_0_LC_8_5_1 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \Lab_UT.didp.curr_LED_0_LC_8_5_1  (
            .in0(N__29724),
            .in1(N__25452),
            .in2(_gnd_net_),
            .in3(N__26152),
            .lcout(\Lab_UT.didp.curr_LEDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29441),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.uu0.counter_gen_label_3__un252_ci_LC_8_5_2 .C_ON=1'b0;
    defparam \resetGen.uu0.counter_gen_label_3__un252_ci_LC_8_5_2 .SEQ_MODE=4'b0000;
    defparam \resetGen.uu0.counter_gen_label_3__un252_ci_LC_8_5_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \resetGen.uu0.counter_gen_label_3__un252_ci_LC_8_5_2  (
            .in0(N__19227),
            .in1(N__19239),
            .in2(_gnd_net_),
            .in3(N__19139),
            .lcout(),
            .ltout(\resetGen.un252_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_3_LC_8_5_3 .C_ON=1'b0;
    defparam \resetGen.reset_count_3_LC_8_5_3 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_3_LC_8_5_3 .LUT_INIT=16'b0100010100010000;
    LogicCell40 \resetGen.reset_count_3_LC_8_5_3  (
            .in0(N__20424),
            .in1(N__19187),
            .in2(N__18940),
            .in3(N__18933),
            .lcout(\resetGen.reset_countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29441),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_1_LC_8_5_4 .C_ON=1'b0;
    defparam \resetGen.reset_count_1_LC_8_5_4 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_1_LC_8_5_4 .LUT_INIT=16'b0000000011000110;
    LogicCell40 \resetGen.reset_count_1_LC_8_5_4  (
            .in0(N__19228),
            .in1(N__19240),
            .in2(N__19192),
            .in3(N__20422),
            .lcout(\resetGen.reset_countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29441),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.uu0.counter_gen_label_2__un241_ci_LC_8_5_5 .C_ON=1'b0;
    defparam \resetGen.uu0.counter_gen_label_2__un241_ci_LC_8_5_5 .SEQ_MODE=4'b0000;
    defparam \resetGen.uu0.counter_gen_label_2__un241_ci_LC_8_5_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \resetGen.uu0.counter_gen_label_2__un241_ci_LC_8_5_5  (
            .in0(N__19238),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19226),
            .lcout(\resetGen.un241_ci ),
            .ltout(\resetGen.un241_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_2_LC_8_5_6 .C_ON=1'b0;
    defparam \resetGen.reset_count_2_LC_8_5_6 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_2_LC_8_5_6 .LUT_INIT=16'b0000000010011100;
    LogicCell40 \resetGen.reset_count_2_LC_8_5_6  (
            .in0(N__19186),
            .in1(N__19140),
            .in2(N__19147),
            .in3(N__20423),
            .lcout(\resetGen.reset_countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29441),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.uu0.delay_line_RNII8EF5_1_LC_8_5_7 .C_ON=1'b0;
    defparam \Lab_UT.uu0.delay_line_RNII8EF5_1_LC_8_5_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.uu0.delay_line_RNII8EF5_1_LC_8_5_7 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \Lab_UT.uu0.delay_line_RNII8EF5_1_LC_8_5_7  (
            .in0(N__19123),
            .in1(N__22146),
            .in2(_gnd_net_),
            .in3(N__23235),
            .lcout(\Lab_UT.uu0.un11_l_count_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_93_LC_8_6_0 .C_ON=1'b0;
    defparam \uu2.bitmap_93_LC_8_6_0 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_93_LC_8_6_0 .LUT_INIT=16'b1111101011110000;
    LogicCell40 \uu2.bitmap_93_LC_8_6_0  (
            .in0(N__19563),
            .in1(_gnd_net_),
            .in2(N__19887),
            .in3(N__19075),
            .lcout(\uu2.bitmapZ0Z_93 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_93C_net ),
            .ce(),
            .sr(N__26048));
    defparam \Lab_UT.didp.Sones_alarm.q_RNIOCVC5_1_LC_8_6_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.Sones_alarm.q_RNIOCVC5_1_LC_8_6_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Sones_alarm.q_RNIOCVC5_1_LC_8_6_1 .LUT_INIT=16'b0101111010110101;
    LogicCell40 \Lab_UT.didp.Sones_alarm.q_RNIOCVC5_1_LC_8_6_1  (
            .in0(N__19354),
            .in1(N__19304),
            .in2(N__19738),
            .in3(N__19265),
            .lcout(\Lab_UT.L3_segment1_1_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Sones_alarm.q_RNIOCVC5_1_1_LC_8_6_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.Sones_alarm.q_RNIOCVC5_1_1_LC_8_6_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Sones_alarm.q_RNIOCVC5_1_1_LC_8_6_2 .LUT_INIT=16'b0100000010000110;
    LogicCell40 \Lab_UT.didp.Sones_alarm.q_RNIOCVC5_1_1_LC_8_6_2  (
            .in0(N__19264),
            .in1(N__19355),
            .in2(N__19316),
            .in3(N__19726),
            .lcout(),
            .ltout(\Lab_UT.L3_segment1_0_i_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_58_LC_8_6_3 .C_ON=1'b0;
    defparam \uu2.bitmap_58_LC_8_6_3 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_58_LC_8_6_3 .LUT_INIT=16'b1100111111001100;
    LogicCell40 \uu2.bitmap_58_LC_8_6_3  (
            .in0(_gnd_net_),
            .in1(N__19851),
            .in2(N__19087),
            .in3(N__19562),
            .lcout(\uu2.bitmapZ0Z_58 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_93C_net ),
            .ce(),
            .sr(N__26048));
    defparam \Lab_UT.didp.Sones_alarm.q_RNIOCVC5_2_1_LC_8_6_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.Sones_alarm.q_RNIOCVC5_2_1_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Sones_alarm.q_RNIOCVC5_2_1_LC_8_6_4 .LUT_INIT=16'b0001110111010111;
    LogicCell40 \Lab_UT.didp.Sones_alarm.q_RNIOCVC5_2_1_LC_8_6_4  (
            .in0(N__19263),
            .in1(N__19353),
            .in2(N__19315),
            .in3(N__19722),
            .lcout(\Lab_UT.L3_segment1_0_i_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Sones_alarm.q_RNIOCVC5_0_1_LC_8_6_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.Sones_alarm.q_RNIOCVC5_0_1_LC_8_6_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Sones_alarm.q_RNIOCVC5_0_1_LC_8_6_5 .LUT_INIT=16'b0011101111101111;
    LogicCell40 \Lab_UT.didp.Sones_alarm.q_RNIOCVC5_0_1_LC_8_6_5  (
            .in0(N__19356),
            .in1(N__19305),
            .in2(N__19739),
            .in3(N__19266),
            .lcout(),
            .ltout(\Lab_UT.L3_segment1_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_221_LC_8_6_6 .C_ON=1'b0;
    defparam \uu2.bitmap_221_LC_8_6_6 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_221_LC_8_6_6 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \uu2.bitmap_221_LC_8_6_6  (
            .in0(N__19561),
            .in1(_gnd_net_),
            .in2(N__19522),
            .in3(N__19857),
            .lcout(\uu2.bitmapZ0Z_221 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_93C_net ),
            .ce(),
            .sr(N__26048));
    defparam \uu2.bitmap_RNI1D952_93_LC_8_6_7 .C_ON=1'b0;
    defparam \uu2.bitmap_RNI1D952_93_LC_8_6_7 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNI1D952_93_LC_8_6_7 .LUT_INIT=16'b1110001000110011;
    LogicCell40 \uu2.bitmap_RNI1D952_93_LC_8_6_7  (
            .in0(N__19519),
            .in1(N__19513),
            .in2(N__19507),
            .in3(N__19491),
            .lcout(\uu2.bitmap_RNI1D952Z0Z_93 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.dicLdAStens_LC_8_7_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.dicLdAStens_LC_8_7_0 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.dictrl.dicLdAStens_LC_8_7_0 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \Lab_UT.dictrl.dicLdAStens_LC_8_7_0  (
            .in0(N__20515),
            .in1(N__20457),
            .in2(N__20476),
            .in3(N__20569),
            .lcout(\Lab_UT.dictrl.dicLdAStensZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29426),
            .ce(),
            .sr(N__23899));
    defparam \Lab_UT.didp.Sones_alarm.q_RNI3O7B1_0_LC_8_7_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.Sones_alarm.q_RNI3O7B1_0_LC_8_7_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Sones_alarm.q_RNI3O7B1_0_LC_8_7_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Lab_UT.didp.Sones_alarm.q_RNI3O7B1_0_LC_8_7_1  (
            .in0(N__29820),
            .in1(N__23075),
            .in2(_gnd_net_),
            .in3(N__19666),
            .lcout(\Lab_UT.Sone_at_0 ),
            .ltout(\Lab_UT.Sone_at_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.segmentUQ_i_a3_0_4_LC_8_7_2 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.segmentUQ_i_a3_0_4_LC_8_7_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.segmentUQ_i_a3_0_4_LC_8_7_2 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \Lab_UT.bcd2segment1.segmentUQ_i_a3_0_4_LC_8_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19330),
            .in3(N__19306),
            .lcout(\Lab_UT.N_77_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Sones_alarm.q_RNI9U7B1_3_LC_8_7_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.Sones_alarm.q_RNI9U7B1_3_LC_8_7_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Sones_alarm.q_RNI9U7B1_3_LC_8_7_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Lab_UT.didp.Sones_alarm.q_RNI9U7B1_3_LC_8_7_3  (
            .in0(N__26188),
            .in1(N__22925),
            .in2(_gnd_net_),
            .in3(N__19669),
            .lcout(\Lab_UT.Sone_at_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Sones_alarm.q_RNI7S7B1_2_LC_8_7_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.Sones_alarm.q_RNI7S7B1_2_LC_8_7_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Sones_alarm.q_RNI7S7B1_2_LC_8_7_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.didp.Sones_alarm.q_RNI7S7B1_2_LC_8_7_4  (
            .in0(N__19667),
            .in1(N__26229),
            .in2(_gnd_net_),
            .in3(N__23036),
            .lcout(\Lab_UT.Sone_at_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Stens_alarm.q_RNIHF5B1_2_LC_8_7_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.Stens_alarm.q_RNIHF5B1_2_LC_8_7_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Stens_alarm.q_RNIHF5B1_2_LC_8_7_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \Lab_UT.didp.Stens_alarm.q_RNIHF5B1_2_LC_8_7_5  (
            .in0(N__25625),
            .in1(N__27162),
            .in2(_gnd_net_),
            .in3(N__19670),
            .lcout(\Lab_UT.Sten_at_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Stens_alarm.q_RNIDB5B1_0_LC_8_7_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.Stens_alarm.q_RNIDB5B1_0_LC_8_7_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Stens_alarm.q_RNIDB5B1_0_LC_8_7_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.didp.Stens_alarm.q_RNIDB5B1_0_LC_8_7_6  (
            .in0(N__19668),
            .in1(N__29689),
            .in2(_gnd_net_),
            .in3(N__25724),
            .lcout(\Lab_UT.Sten_at_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Stens_alarm.q_RNIJH5B1_3_LC_8_7_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.Stens_alarm.q_RNIJH5B1_3_LC_8_7_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Stens_alarm.q_RNIJH5B1_3_LC_8_7_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Lab_UT.didp.Stens_alarm.q_RNIJH5B1_3_LC_8_7_7  (
            .in0(N__27126),
            .in1(N__22979),
            .in2(_gnd_net_),
            .in3(N__19671),
            .lcout(\Lab_UT.Sten_at_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Stens_alarm.q_RNIFD5B1_1_LC_8_8_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.Stens_alarm.q_RNIFD5B1_1_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Stens_alarm.q_RNIFD5B1_1_LC_8_8_0 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \Lab_UT.didp.Stens_alarm.q_RNIFD5B1_1_LC_8_8_0  (
            .in0(N__19660),
            .in1(_gnd_net_),
            .in2(N__25809),
            .in3(N__27872),
            .lcout(\Lab_UT.Sten_at_1 ),
            .ltout(\Lab_UT.Sten_at_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment2.segmentUQ_0_5_LC_8_8_1 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment2.segmentUQ_0_5_LC_8_8_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment2.segmentUQ_0_5_LC_8_8_1 .LUT_INIT=16'b0010100000110010;
    LogicCell40 \Lab_UT.bcd2segment2.segmentUQ_0_5_LC_8_8_1  (
            .in0(N__20030),
            .in1(N__19987),
            .in2(N__19954),
            .in3(N__19923),
            .lcout(\Lab_UT.segmentUQ_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_0_ret_11_RNIA2D93_LC_8_8_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_11_RNIA2D93_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_0_ret_11_RNIA2D93_LC_8_8_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_11_RNIA2D93_LC_8_8_4  (
            .in0(N__20824),
            .in1(N__27811),
            .in2(_gnd_net_),
            .in3(N__27300),
            .lcout(\Lab_UT.dicLdStens_latmux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_0_ret_14_RNID3D61_LC_8_8_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_14_RNID3D61_LC_8_8_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_0_ret_14_RNID3D61_LC_8_8_5 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_14_RNID3D61_LC_8_8_5  (
            .in0(N__26675),
            .in1(N__24172),
            .in2(N__29491),
            .in3(N__23646),
            .lcout(\Lab_UT.dictrl.L3_segment1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Sones_alarm.q_RNI5Q7B1_1_LC_8_8_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.Sones_alarm.q_RNI5Q7B1_1_LC_8_8_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Sones_alarm.q_RNI5Q7B1_1_LC_8_8_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \Lab_UT.didp.Sones_alarm.q_RNI5Q7B1_1_LC_8_8_7  (
            .in0(N__23059),
            .in1(N__28104),
            .in2(_gnd_net_),
            .in3(N__19659),
            .lcout(\Lab_UT.Sone_at_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_0_ret_3_RNI9MVL_0_LC_8_9_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_3_RNI9MVL_0_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_0_ret_3_RNI9MVL_0_LC_8_9_0 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_3_RNI9MVL_0_LC_8_9_0  (
            .in0(N__26676),
            .in1(N__23476),
            .in2(_gnd_net_),
            .in3(N__23161),
            .lcout(\Lab_UT.dictrl.r_enable1_2_i_m ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.r_alarm_or_time_RNI9J3I_LC_8_9_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.r_alarm_or_time_RNI9J3I_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.r_alarm_or_time_RNI9J3I_LC_8_9_1 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \Lab_UT.dictrl.r_alarm_or_time_RNI9J3I_LC_8_9_1  (
            .in0(N__24157),
            .in1(N__23637),
            .in2(_gnd_net_),
            .in3(N__20223),
            .lcout(\Lab_UT.alarm_or_time_0 ),
            .ltout(\Lab_UT.alarm_or_time_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Mtens_alarm.q_RNI5TK11_2_LC_8_9_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mtens_alarm.q_RNI5TK11_2_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Mtens_alarm.q_RNI5TK11_2_LC_8_9_2 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \Lab_UT.didp.Mtens_alarm.q_RNI5TK11_2_LC_8_9_2  (
            .in0(N__25844),
            .in1(_gnd_net_),
            .in2(N__19612),
            .in3(N__26873),
            .lcout(\Lab_UT.Mten_at_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.dicLdStens_LC_8_9_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.dicLdStens_LC_8_9_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.dicLdStens_LC_8_9_3 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \Lab_UT.dictrl.dicLdStens_LC_8_9_3  (
            .in0(N__29939),
            .in1(N__23092),
            .in2(N__23113),
            .in3(N__29882),
            .lcout(\Lab_UT.dicLdStens ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29409),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_0_ret_3_RNI9MVL_LC_8_9_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_3_RNI9MVL_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_0_ret_3_RNI9MVL_LC_8_9_4 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_3_RNI9MVL_LC_8_9_4  (
            .in0(N__26677),
            .in1(N__23477),
            .in2(_gnd_net_),
            .in3(N__23162),
            .lcout(\Lab_UT.dictrl.r_enable1_2_m ),
            .ltout(\Lab_UT.dictrl.r_enable1_2_m_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.r_enable2_LC_8_9_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.r_enable2_LC_8_9_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.r_enable2_LC_8_9_5 .LUT_INIT=16'b1111101101010001;
    LogicCell40 \Lab_UT.dictrl.r_enable2_LC_8_9_5  (
            .in0(N__23440),
            .in1(N__20260),
            .in2(N__20191),
            .in3(N__20179),
            .lcout(\Lab_UT.dictrl.r_enableZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29409),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_0_ret_29_RNIPGJ2_LC_8_9_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_29_RNIPGJ2_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_0_ret_29_RNIPGJ2_LC_8_9_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_29_RNIPGJ2_LC_8_9_6  (
            .in0(_gnd_net_),
            .in1(N__23439),
            .in2(_gnd_net_),
            .in3(N__26149),
            .lcout(\Lab_UT.dictrl.g0_i_a4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.r_enable2_RNI8DR61_LC_8_9_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.r_enable2_RNI8DR61_LC_8_9_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.r_enable2_RNI8DR61_LC_8_9_7 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \Lab_UT.dictrl.r_enable2_RNI8DR61_LC_8_9_7  (
            .in0(N__24158),
            .in1(N__20178),
            .in2(N__23170),
            .in3(N__23638),
            .lcout(\Lab_UT.dictrl.enableSeg2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_0_ret_22_LC_8_10_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_22_LC_8_10_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.currState_0_ret_22_LC_8_10_0 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_22_LC_8_10_0  (
            .in0(N__20125),
            .in1(N__24687),
            .in2(_gnd_net_),
            .in3(N__20119),
            .lcout(\Lab_UT.un1_r_Sone_init5_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29402),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_ret_0_LC_8_10_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_ret_0_LC_8_10_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.currState_ret_0_LC_8_10_1 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \Lab_UT.dictrl.currState_ret_0_LC_8_10_1  (
            .in0(N__24686),
            .in1(N__20767),
            .in2(N__24730),
            .in3(N__21606),
            .lcout(\Lab_UT.dictrl.r_dicLdMtens19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29402),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_0_ret_23_LC_8_10_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_23_LC_8_10_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.currState_0_ret_23_LC_8_10_2 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_23_LC_8_10_2  (
            .in0(N__20561),
            .in1(N__24726),
            .in2(_gnd_net_),
            .in3(N__24688),
            .lcout(\Lab_UT.dictrl.r_dicLdMtens23_i_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29402),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.r_enable2_RNO_1_LC_8_10_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.r_enable2_RNO_1_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.r_enable2_RNO_1_LC_8_10_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Lab_UT.dictrl.r_enable2_RNO_1_LC_8_10_3  (
            .in0(N__20086),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20206),
            .lcout(),
            .ltout(\Lab_UT.dictrl.r_enable2_3_iv_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.r_enable2_RNO_0_LC_8_10_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.r_enable2_RNO_0_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.r_enable2_RNO_0_LC_8_10_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.r_enable2_RNO_0_LC_8_10_4  (
            .in0(N__20212),
            .in1(N__20235),
            .in2(N__20263),
            .in3(N__23595),
            .lcout(\Lab_UT.dictrl.r_enable2_3_iv_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.r_alarm_or_time_RNO_0_LC_8_10_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.r_alarm_or_time_RNO_0_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.r_alarm_or_time_RNO_0_LC_8_10_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.dictrl.r_alarm_or_time_RNO_0_LC_8_10_6  (
            .in0(_gnd_net_),
            .in1(N__20251),
            .in2(_gnd_net_),
            .in3(N__20236),
            .lcout(),
            .ltout(\Lab_UT.dictrl.un1_r_dicLdMtens19_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.r_alarm_or_time_LC_8_10_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.r_alarm_or_time_LC_8_10_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.r_alarm_or_time_LC_8_10_7 .LUT_INIT=16'b0100010100000001;
    LogicCell40 \Lab_UT.dictrl.r_alarm_or_time_LC_8_10_7  (
            .in0(N__23478),
            .in1(N__23435),
            .in2(N__20227),
            .in3(N__20224),
            .lcout(\Lab_UT.dictrl.r_alarm_or_timeZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29402),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_0_ret_12_LC_8_11_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_12_LC_8_11_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.currState_0_ret_12_LC_8_11_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_12_LC_8_11_0  (
            .in0(N__21615),
            .in1(N__20661),
            .in2(N__20806),
            .in3(N__21095),
            .lcout(\Lab_UT.dictrl.r_dicLdMtens15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29396),
            .ce(),
            .sr(N__26071));
    defparam \Lab_UT.dictrl.currState_0_ret_16_LC_8_11_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_16_LC_8_11_1 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.currState_0_ret_16_LC_8_11_1 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_16_LC_8_11_1  (
            .in0(N__21091),
            .in1(N__21619),
            .in2(N__20810),
            .in3(N__20665),
            .lcout(\Lab_UT.dictrl.r_dicLdMtens18_i_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29396),
            .ce(),
            .sr(N__26071));
    defparam \Lab_UT.dictrl.currState_0_ret_18_LC_8_11_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_18_LC_8_11_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.currState_0_ret_18_LC_8_11_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_18_LC_8_11_2  (
            .in0(N__21616),
            .in1(N__20662),
            .in2(N__20807),
            .in3(N__21096),
            .lcout(\Lab_UT.dictrl.r_dicLdMtens17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29396),
            .ce(),
            .sr(N__26071));
    defparam \Lab_UT.dictrl.currState_0_ret_19_LC_8_11_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_19_LC_8_11_3 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.currState_0_ret_19_LC_8_11_3 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_19_LC_8_11_3  (
            .in0(N__21092),
            .in1(N__21620),
            .in2(N__20811),
            .in3(N__20666),
            .lcout(\Lab_UT.dictrl.r_dicLdMtens17_i_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29396),
            .ce(),
            .sr(N__26071));
    defparam \Lab_UT.dictrl.currState_0_ret_6_LC_8_11_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_6_LC_8_11_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.currState_0_ret_6_LC_8_11_4 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_6_LC_8_11_4  (
            .in0(N__21617),
            .in1(N__20663),
            .in2(N__20808),
            .in3(N__21097),
            .lcout(\Lab_UT.dictrl.r_dicLdMtens14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29396),
            .ce(),
            .sr(N__26071));
    defparam \Lab_UT.dictrl.currState_0_ret_7_LC_8_11_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_7_LC_8_11_5 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.currState_0_ret_7_LC_8_11_5 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_7_LC_8_11_5  (
            .in0(N__21093),
            .in1(N__21621),
            .in2(N__20812),
            .in3(N__20667),
            .lcout(\Lab_UT.dictrl.r_dicLdMtens14_i_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29396),
            .ce(),
            .sr(N__26071));
    defparam \Lab_UT.dictrl.currState_0_ret_11_LC_8_11_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_11_LC_8_11_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.currState_0_ret_11_LC_8_11_6 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_11_LC_8_11_6  (
            .in0(N__21614),
            .in1(N__20660),
            .in2(N__20805),
            .in3(N__21094),
            .lcout(\Lab_UT.dictrl.r_dicLdMtens16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29396),
            .ce(),
            .sr(N__26071));
    defparam \Lab_UT.dictrl.currState_0_ret_15_LC_8_11_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_15_LC_8_11_7 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.currState_0_ret_15_LC_8_11_7 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_15_LC_8_11_7  (
            .in0(N__21090),
            .in1(N__21618),
            .in2(N__20809),
            .in3(N__20664),
            .lcout(\Lab_UT.dictrl.un2_dicAlarmTrig_i_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29396),
            .ce(),
            .sr(N__26071));
    defparam \Lab_UT.dictrl.currState_0_ret_18_RNIH2D93_LC_8_12_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_18_RNIH2D93_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_0_ret_18_RNIH2D93_LC_8_12_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_18_RNIH2D93_LC_8_12_0  (
            .in0(N__20578),
            .in1(N__27806),
            .in2(_gnd_net_),
            .in3(N__27559),
            .lcout(\Lab_UT.dicLdSones_latmux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.dicLdAMones_LC_8_12_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.dicLdAMones_LC_8_12_1 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.dictrl.dicLdAMones_LC_8_12_1 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \Lab_UT.dictrl.dicLdAMones_LC_8_12_1  (
            .in0(N__20562),
            .in1(N__20530),
            .in2(N__20539),
            .in3(N__20518),
            .lcout(\Lab_UT.dictrl.dicLdAMonesZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29392),
            .ce(),
            .sr(N__23920));
    defparam \Lab_UT.dictrl.currState_ret_7_RNIUEJQ4_LC_8_12_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_ret_7_RNIUEJQ4_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_ret_7_RNIUEJQ4_LC_8_12_2 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \Lab_UT.dictrl.currState_ret_7_RNIUEJQ4_LC_8_12_2  (
            .in0(N__23913),
            .in1(N__27807),
            .in2(_gnd_net_),
            .in3(N__27560),
            .lcout(\Lab_UT.dictrl.dicLdAMones_rst ),
            .ltout(\Lab_UT.dictrl.dicLdAMones_rst_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.dicLdAMones_RNI3BNL5_LC_8_12_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.dicLdAMones_RNI3BNL5_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.dicLdAMones_RNI3BNL5_LC_8_12_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \Lab_UT.dictrl.dicLdAMones_RNI3BNL5_LC_8_12_3  (
            .in0(_gnd_net_),
            .in1(N__20529),
            .in2(N__20521),
            .in3(N__20517),
            .lcout(\Lab_UT.ld_enable_AMones ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.dicLdAStens_RNI7OAH5_LC_8_12_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.dicLdAStens_RNI7OAH5_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.dicLdAStens_RNI7OAH5_LC_8_12_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Lab_UT.dictrl.dicLdAStens_RNI7OAH5_LC_8_12_4  (
            .in0(N__20516),
            .in1(N__20475),
            .in2(_gnd_net_),
            .in3(N__20458),
            .lcout(\Lab_UT.ld_enable_AStens ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.escKey_LC_8_12_5 .C_ON=1'b0;
    defparam \resetGen.escKey_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \resetGen.escKey_LC_8_12_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \resetGen.escKey_LC_8_12_5  (
            .in0(N__27808),
            .in1(N__21118),
            .in2(_gnd_net_),
            .in3(N__25435),
            .lcout(\resetGen.escKeyZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__m5_LC_8_12_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__m5_LC_8_12_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__m5_LC_8_12_6 .LUT_INIT=16'b1011101101010101;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__m5_LC_8_12_6  (
            .in0(N__20395),
            .in1(N__24476),
            .in2(_gnd_net_),
            .in3(N__20299),
            .lcout(\Lab_UT.dictrl.N_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.r_enable3_RNO_0_LC_8_12_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.r_enable3_RNO_0_LC_8_12_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.r_enable3_RNO_0_LC_8_12_7 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \Lab_UT.dictrl.r_enable3_RNO_0_LC_8_12_7  (
            .in0(N__21325),
            .in1(N__21319),
            .in2(_gnd_net_),
            .in3(N__23686),
            .lcout(\Lab_UT.dictrl.r_enable3_3_iv_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_RNI86KI_6_LC_8_13_0 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_RNI86KI_6_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.shifter_RNI86KI_6_LC_8_13_0 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \buart.Z_rx.shifter_RNI86KI_6_LC_8_13_0  (
            .in0(_gnd_net_),
            .in1(N__24295),
            .in2(_gnd_net_),
            .in3(N__28508),
            .lcout(),
            .ltout(\buart.Z_rx.G_30_0_o3_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_RNIV4BN3_7_LC_8_13_1 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_RNIV4BN3_7_LC_8_13_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.shifter_RNIV4BN3_7_LC_8_13_1 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \buart.Z_rx.shifter_RNIV4BN3_7_LC_8_13_1  (
            .in0(N__21634),
            .in1(N__25395),
            .in2(N__21295),
            .in3(N__21292),
            .lcout(),
            .ltout(N_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_0_ret_21_RNI88818_LC_8_13_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_21_RNI88818_LC_8_13_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_0_ret_21_RNI88818_LC_8_13_2 .LUT_INIT=16'b1000000010001111;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_21_RNI88818_LC_8_13_2  (
            .in0(N__21260),
            .in1(N__24475),
            .in2(N__21136),
            .in3(N__24011),
            .lcout(\Lab_UT.dictrl.N_21_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.escKey_4_LC_8_13_3 .C_ON=1'b0;
    defparam \resetGen.escKey_4_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \resetGen.escKey_4_LC_8_13_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \resetGen.escKey_4_LC_8_13_3  (
            .in0(N__28509),
            .in1(N__24447),
            .in2(N__24310),
            .in3(N__25396),
            .lcout(\resetGen.escKey_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_0_rep2_LC_8_13_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_0_rep2_LC_8_13_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.currState_2_0_rep2_LC_8_13_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Lab_UT.dictrl.currState_2_0_rep2_LC_8_13_4  (
            .in0(_gnd_net_),
            .in1(N__24695),
            .in2(_gnd_net_),
            .in3(N__21107),
            .lcout(\Lab_UT.dictrl.currState_0_rep2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29386),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_14_LC_8_13_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_14_LC_8_13_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_14_LC_8_13_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__g0_14_LC_8_13_6  (
            .in0(N__28743),
            .in1(N__28507),
            .in2(N__28947),
            .in3(N__25304),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_7_LC_8_13_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_7_LC_8_13_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g0_7_LC_8_13_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__g0_7_LC_8_13_7  (
            .in0(N__24296),
            .in1(N__20900),
            .in2(N__20860),
            .in3(N__24890),
            .lcout(\Lab_UT.dictrl.g0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.decoder.de_littleL_4_LC_8_14_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.decoder.de_littleL_4_LC_8_14_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.decoder.de_littleL_4_LC_8_14_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Lab_UT.dictrl.decoder.de_littleL_4_LC_8_14_0  (
            .in0(N__21442),
            .in1(N__21346),
            .in2(N__21831),
            .in3(N__20838),
            .lcout(\Lab_UT.dictrl.de_littleL_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__g1_6_LC_8_14_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g1_6_LC_8_14_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g1_6_LC_8_14_1 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__g1_6_LC_8_14_1  (
            .in0(N__21347),
            .in1(N__21443),
            .in2(N__21781),
            .in3(N__21819),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g1_5_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__g1_2_LC_8_14_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g1_2_LC_8_14_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g1_2_LC_8_14_2 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__g1_2_LC_8_14_2  (
            .in0(N__21407),
            .in1(N__21649),
            .in2(N__21718),
            .in3(N__24308),
            .lcout(\Lab_UT.dictrl.g1_7_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_1_3_0__g1_3_LC_8_14_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g1_3_LC_8_14_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_1_3_0__g1_3_LC_8_14_3 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \Lab_UT.dictrl.nextState_1_3_0__g1_3_LC_8_14_3  (
            .in0(N__21640),
            .in1(N__21699),
            .in2(_gnd_net_),
            .in3(N__21924),
            .lcout(\Lab_UT.dictrl.g1_4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_3_fast_3_LC_8_14_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_3_fast_3_LC_8_14_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.currState_3_fast_3_LC_8_14_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.dictrl.currState_3_fast_3_LC_8_14_4  (
            .in0(_gnd_net_),
            .in1(N__24704),
            .in2(_gnd_net_),
            .in3(N__21623),
            .lcout(\Lab_UT.dictrl.currState_fast_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29382),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_RNID9851_4_LC_8_14_5 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_RNID9851_4_LC_8_14_5 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.shifter_RNID9851_4_LC_8_14_5 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \buart.Z_rx.shifter_RNID9851_4_LC_8_14_5  (
            .in0(N__24443),
            .in1(N__28753),
            .in2(N__28964),
            .in3(N__25303),
            .lcout(\buart.Z_rx.G_30_0_o3_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_3_3_LC_8_14_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_3_3_LC_8_14_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.currState_3_3_LC_8_14_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.dictrl.currState_3_3_LC_8_14_6  (
            .in0(_gnd_net_),
            .in1(N__24703),
            .in2(_gnd_net_),
            .in3(N__21622),
            .lcout(\Lab_UT.dictrl.currStateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29382),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.decoder.g0_12_LC_8_14_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.decoder.g0_12_LC_8_14_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.decoder.g0_12_LC_8_14_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Lab_UT.dictrl.decoder.g0_12_LC_8_14_7  (
            .in0(N__21445),
            .in1(N__21925),
            .in2(N__21987),
            .in3(N__21406),
            .lcout(\Lab_UT.dictrl.decoder.g0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_0_LC_8_15_0 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_LC_8_15_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_0_LC_8_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_0_LC_8_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28771),
            .lcout(bu_rx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29378),
            .ce(N__25424),
            .sr(N__26101));
    defparam \buart.Z_rx.shifter_0_rep1_LC_8_15_2 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_rep1_LC_8_15_2 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_0_rep1_LC_8_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_0_rep1_LC_8_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28772),
            .lcout(bu_rx_data_0_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29378),
            .ce(N__25424),
            .sr(N__26101));
    defparam \buart.Z_rx.shifter_6_rep1_LC_8_15_3 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_6_rep1_LC_8_15_3 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_6_rep1_LC_8_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_6_rep1_LC_8_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25377),
            .lcout(bu_rx_data_6_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29378),
            .ce(N__25424),
            .sr(N__26101));
    defparam \buart.Z_rx.shifter_3_LC_8_15_4 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_3_LC_8_15_4 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_3_LC_8_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_3_LC_8_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25301),
            .lcout(bu_rx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29378),
            .ce(N__25424),
            .sr(N__26101));
    defparam \buart.Z_rx.shifter_5_rep1_LC_8_15_5 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_5_rep1_LC_8_15_5 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_5_rep1_LC_8_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_5_rep1_LC_8_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24300),
            .lcout(bu_rx_data_5_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29378),
            .ce(N__25424),
            .sr(N__26101));
    defparam \buart.Z_rx.shifter_fast_3_LC_8_15_6 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_3_LC_8_15_6 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_fast_3_LC_8_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_fast_3_LC_8_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25302),
            .lcout(bu_rx_data_fast_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29378),
            .ce(N__25424),
            .sr(N__26101));
    defparam \buart.Z_rx.shifter_7_rep1_LC_8_15_7 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_7_rep1_LC_8_15_7 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_7_rep1_LC_8_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_7_rep1_LC_8_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21876),
            .lcout(bu_rx_data_7_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29378),
            .ce(N__25424),
            .sr(N__26101));
    defparam \Lab_UT.uu0.l_count_1_LC_9_1_0 .C_ON=1'b0;
    defparam \Lab_UT.uu0.l_count_1_LC_9_1_0 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.uu0.l_count_1_LC_9_1_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \Lab_UT.uu0.l_count_1_LC_9_1_0  (
            .in0(N__22093),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22521),
            .lcout(\Lab_UT.uu0.l_countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29476),
            .ce(N__22171),
            .sr(N__26105));
    defparam \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_1_LC_9_1_1 .C_ON=1'b0;
    defparam \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_1_LC_9_1_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_1_LC_9_1_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_1_LC_9_1_1  (
            .in0(N__22519),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22092),
            .lcout(\Lab_UT.uu0.un44_ci ),
            .ltout(\Lab_UT.uu0.un44_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.uu0.l_count_3_LC_9_1_2 .C_ON=1'b0;
    defparam \Lab_UT.uu0.l_count_3_LC_9_1_2 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.uu0.l_count_3_LC_9_1_2 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \Lab_UT.uu0.l_count_3_LC_9_1_2  (
            .in0(N__22243),
            .in1(N__22260),
            .in2(N__21784),
            .in3(N__23222),
            .lcout(\Lab_UT.uu0.l_countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29476),
            .ce(N__22171),
            .sr(N__26105));
    defparam \Lab_UT.uu0.l_count_0_LC_9_1_4 .C_ON=1'b0;
    defparam \Lab_UT.uu0.l_count_0_LC_9_1_4 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.uu0.l_count_0_LC_9_1_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Lab_UT.uu0.l_count_0_LC_9_1_4  (
            .in0(_gnd_net_),
            .in1(N__22520),
            .in2(_gnd_net_),
            .in3(N__23220),
            .lcout(\Lab_UT.uu0.l_countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29476),
            .ce(N__22171),
            .sr(N__26105));
    defparam \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_9_1_5 .C_ON=1'b0;
    defparam \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_9_1_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_9_1_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_9_1_5  (
            .in0(N__22259),
            .in1(N__22242),
            .in2(N__22522),
            .in3(N__22091),
            .lcout(\Lab_UT.uu0.un66_ci ),
            .ltout(\Lab_UT.uu0.un66_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.uu0.l_count_4_LC_9_1_6 .C_ON=1'b0;
    defparam \Lab_UT.uu0.l_count_4_LC_9_1_6 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.uu0.l_count_4_LC_9_1_6 .LUT_INIT=16'b0000000000111100;
    LogicCell40 \Lab_UT.uu0.l_count_4_LC_9_1_6  (
            .in0(_gnd_net_),
            .in1(N__22215),
            .in2(N__22219),
            .in3(N__23221),
            .lcout(\Lab_UT.uu0.l_countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29476),
            .ce(N__22171),
            .sr(N__26105));
    defparam \Lab_UT.uu0.l_count_5_LC_9_1_7 .C_ON=1'b0;
    defparam \Lab_UT.uu0.l_count_5_LC_9_1_7 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.uu0.l_count_5_LC_9_1_7 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \Lab_UT.uu0.l_count_5_LC_9_1_7  (
            .in0(N__22216),
            .in1(N__22193),
            .in2(_gnd_net_),
            .in3(N__22129),
            .lcout(\Lab_UT.uu0.l_countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29476),
            .ce(N__22171),
            .sr(N__26105));
    defparam \Lab_UT.uu0.delay_line_0_LC_9_2_0 .C_ON=1'b0;
    defparam \Lab_UT.uu0.delay_line_0_LC_9_2_0 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.uu0.delay_line_0_LC_9_2_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.uu0.delay_line_0_LC_9_2_0  (
            .in0(N__22594),
            .in1(N__25210),
            .in2(N__22111),
            .in3(N__22537),
            .lcout(\Lab_UT.uu0.delay_lineZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29472),
            .ce(),
            .sr(N__26104));
    defparam \Lab_UT.uu0.l_precount_3_LC_9_2_1 .C_ON=1'b0;
    defparam \Lab_UT.uu0.l_precount_3_LC_9_2_1 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.uu0.l_precount_3_LC_9_2_1 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \Lab_UT.uu0.l_precount_3_LC_9_2_1  (
            .in0(N__22539),
            .in1(N__22109),
            .in2(N__25216),
            .in3(N__22597),
            .lcout(\Lab_UT.uu0.l_precountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29472),
            .ce(),
            .sr(N__26104));
    defparam \Lab_UT.uu0.l_count_RNIS3Q51_5_LC_9_2_2 .C_ON=1'b0;
    defparam \Lab_UT.uu0.l_count_RNIS3Q51_5_LC_9_2_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.uu0.l_count_RNIS3Q51_5_LC_9_2_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Lab_UT.uu0.l_count_RNIS3Q51_5_LC_9_2_2  (
            .in0(N__22593),
            .in1(N__22127),
            .in2(N__22110),
            .in3(N__22090),
            .lcout(),
            .ltout(\Lab_UT.uu0.un4_l_count_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.uu0.l_count_RNIC7FP1_18_LC_9_2_3 .C_ON=1'b0;
    defparam \Lab_UT.uu0.l_count_RNIC7FP1_18_LC_9_2_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.uu0.l_count_RNIC7FP1_18_LC_9_2_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.uu0.l_count_RNIC7FP1_18_LC_9_2_3  (
            .in0(N__22075),
            .in1(N__22055),
            .in2(N__22039),
            .in3(N__22033),
            .lcout(),
            .ltout(\Lab_UT.uu0.un4_l_count_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.uu0.l_count_RNIRSCC5_3_LC_9_2_4 .C_ON=1'b0;
    defparam \Lab_UT.uu0.l_count_RNIRSCC5_3_LC_9_2_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.uu0.l_count_RNIRSCC5_3_LC_9_2_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.uu0.l_count_RNIRSCC5_3_LC_9_2_4  (
            .in0(N__22498),
            .in1(N__22018),
            .in2(N__22009),
            .in3(N__22006),
            .lcout(\Lab_UT.uu0.un4_l_count_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.uu0.l_precount_1_LC_9_2_5 .C_ON=1'b0;
    defparam \Lab_UT.uu0.l_precount_1_LC_9_2_5 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.uu0.l_precount_1_LC_9_2_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \Lab_UT.uu0.l_precount_1_LC_9_2_5  (
            .in0(N__25211),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22595),
            .lcout(\Lab_UT.uu0.l_precountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29472),
            .ce(),
            .sr(N__26104));
    defparam \Lab_UT.uu0.l_precount_2_LC_9_2_6 .C_ON=1'b0;
    defparam \Lab_UT.uu0.l_precount_2_LC_9_2_6 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.uu0.l_precount_2_LC_9_2_6 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \Lab_UT.uu0.l_precount_2_LC_9_2_6  (
            .in0(N__22596),
            .in1(N__25212),
            .in2(_gnd_net_),
            .in3(N__22538),
            .lcout(\Lab_UT.uu0.l_precountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29472),
            .ce(),
            .sr(N__26104));
    defparam \Lab_UT.uu0.l_count_RNIM5011_11_LC_9_2_7 .C_ON=1'b0;
    defparam \Lab_UT.uu0.l_count_RNIM5011_11_LC_9_2_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.uu0.l_count_RNIM5011_11_LC_9_2_7 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \Lab_UT.uu0.l_count_RNIM5011_11_LC_9_2_7  (
            .in0(N__22576),
            .in1(N__22556),
            .in2(N__22540),
            .in3(N__22515),
            .lcout(\Lab_UT.uu0.un4_l_count_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_5_LC_9_3_0 .C_ON=1'b0;
    defparam \uu2.w_addr_user_5_LC_9_3_0 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_5_LC_9_3_0 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.w_addr_user_5_LC_9_3_0  (
            .in0(N__22428),
            .in1(N__22396),
            .in2(N__22462),
            .in3(N__22486),
            .lcout(\uu2.w_addr_userZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_5C_net ),
            .ce(),
            .sr(N__22326));
    defparam \uu2.w_addr_user_4_LC_9_3_1 .C_ON=1'b0;
    defparam \uu2.w_addr_user_4_LC_9_3_1 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_4_LC_9_3_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \uu2.w_addr_user_4_LC_9_3_1  (
            .in0(N__22395),
            .in1(N__22455),
            .in2(_gnd_net_),
            .in3(N__22427),
            .lcout(\uu2.w_addr_userZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_5C_net ),
            .ce(),
            .sr(N__22326));
    defparam \uu2.w_addr_user_6_LC_9_3_2 .C_ON=1'b0;
    defparam \uu2.w_addr_user_6_LC_9_3_2 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_6_LC_9_3_2 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.w_addr_user_6_LC_9_3_2  (
            .in0(N__22429),
            .in1(N__22397),
            .in2(N__22378),
            .in3(N__22350),
            .lcout(\uu2.w_addr_userZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_5C_net ),
            .ce(),
            .sr(N__22326));
    defparam \Lab_UT.display.cnt_RNIFA8M_0_2_LC_9_4_0 .C_ON=1'b0;
    defparam \Lab_UT.display.cnt_RNIFA8M_0_2_LC_9_4_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.display.cnt_RNIFA8M_0_2_LC_9_4_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.display.cnt_RNIFA8M_0_2_LC_9_4_0  (
            .in0(_gnd_net_),
            .in1(N__26511),
            .in2(_gnd_net_),
            .in3(N__26426),
            .lcout(\Lab_UT.display.N_150 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.display.rdy_LC_9_4_1 .C_ON=1'b0;
    defparam \Lab_UT.display.rdy_LC_9_4_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.display.rdy_LC_9_4_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Lab_UT.display.rdy_LC_9_4_1  (
            .in0(N__26428),
            .in1(N__26337),
            .in2(N__26515),
            .in3(N__26734),
            .lcout(L3_tx_data_rdy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29457),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.display.dOut_6_LC_9_4_2 .C_ON=1'b0;
    defparam \Lab_UT.display.dOut_6_LC_9_4_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.display.dOut_6_LC_9_4_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \Lab_UT.display.dOut_6_LC_9_4_2  (
            .in0(N__27424),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22854),
            .lcout(L3_tx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29457),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.display.cnt_RNI5EC11_0_LC_9_4_3 .C_ON=1'b0;
    defparam \Lab_UT.display.cnt_RNI5EC11_0_LC_9_4_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.display.cnt_RNI5EC11_0_LC_9_4_3 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \Lab_UT.display.cnt_RNI5EC11_0_LC_9_4_3  (
            .in0(_gnd_net_),
            .in1(N__25565),
            .in2(_gnd_net_),
            .in3(N__26335),
            .lcout(\Lab_UT.display.N_88 ),
            .ltout(\Lab_UT.display.N_88_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.display.dOut_1_LC_9_4_4 .C_ON=1'b0;
    defparam \Lab_UT.display.dOut_1_LC_9_4_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.display.dOut_1_LC_9_4_4 .LUT_INIT=16'b1111111111001110;
    LogicCell40 \Lab_UT.display.dOut_1_LC_9_4_4  (
            .in0(N__23131),
            .in1(N__25753),
            .in2(N__22669),
            .in3(N__22888),
            .lcout(L3_tx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29457),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.display.dOut_RNO_0_4_LC_9_4_5 .C_ON=1'b0;
    defparam \Lab_UT.display.dOut_RNO_0_4_LC_9_4_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.display.dOut_RNO_0_4_LC_9_4_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.display.dOut_RNO_0_4_LC_9_4_5  (
            .in0(_gnd_net_),
            .in1(N__27367),
            .in2(_gnd_net_),
            .in3(N__25566),
            .lcout(),
            .ltout(\Lab_UT.display.N_120_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.display.dOut_4_LC_9_4_6 .C_ON=1'b0;
    defparam \Lab_UT.display.dOut_4_LC_9_4_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.display.dOut_4_LC_9_4_6 .LUT_INIT=16'b0000000100000011;
    LogicCell40 \Lab_UT.display.dOut_4_LC_9_4_6  (
            .in0(N__26336),
            .in1(N__25551),
            .in2(N__22642),
            .in3(N__26427),
            .lcout(L3_tx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29457),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.display.dOut_5_LC_9_4_7 .C_ON=1'b0;
    defparam \Lab_UT.display.dOut_5_LC_9_4_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.display.dOut_5_LC_9_4_7 .LUT_INIT=16'b0001010100010001;
    LogicCell40 \Lab_UT.display.dOut_5_LC_9_4_7  (
            .in0(N__25552),
            .in1(N__25567),
            .in2(N__26341),
            .in3(N__23614),
            .lcout(L3_tx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29457),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.display.dOut_RNO_1_2_LC_9_5_0 .C_ON=1'b0;
    defparam \Lab_UT.display.dOut_RNO_1_2_LC_9_5_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.display.dOut_RNO_1_2_LC_9_5_0 .LUT_INIT=16'b0010001011110010;
    LogicCell40 \Lab_UT.display.dOut_RNO_1_2_LC_9_5_0  (
            .in0(N__26542),
            .in1(N__22733),
            .in2(N__22881),
            .in3(N__23037),
            .lcout(\Lab_UT.display.dOutP_0_iv_i_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.display.dOut_RNO_1_0_LC_9_5_1 .C_ON=1'b0;
    defparam \Lab_UT.display.dOut_RNO_1_0_LC_9_5_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.display.dOut_RNO_1_0_LC_9_5_1 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \Lab_UT.display.dOut_RNO_1_0_LC_9_5_1  (
            .in0(N__26541),
            .in1(N__22874),
            .in2(N__22764),
            .in3(N__23076),
            .lcout(\Lab_UT.display.dOutP_0_iv_i_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.display.cnt_RNIFA8M_1_2_LC_9_5_2 .C_ON=1'b0;
    defparam \Lab_UT.display.cnt_RNIFA8M_1_2_LC_9_5_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.display.cnt_RNIFA8M_1_2_LC_9_5_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Lab_UT.display.cnt_RNIFA8M_1_2_LC_9_5_2  (
            .in0(_gnd_net_),
            .in1(N__26509),
            .in2(_gnd_net_),
            .in3(N__26425),
            .lcout(\Lab_UT.display.N_153 ),
            .ltout(\Lab_UT.display.N_153_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.display.dOut_RNO_1_3_LC_9_5_3 .C_ON=1'b0;
    defparam \Lab_UT.display.dOut_RNO_1_3_LC_9_5_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.display.dOut_RNO_1_3_LC_9_5_3 .LUT_INIT=16'b1101110011001100;
    LogicCell40 \Lab_UT.display.dOut_RNO_1_3_LC_9_5_3  (
            .in0(N__22984),
            .in1(N__25504),
            .in2(N__22600),
            .in3(N__26332),
            .lcout(\Lab_UT.display.dOutP_0_iv_i_2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.display.dOut_RNO_1_1_LC_9_5_4 .C_ON=1'b0;
    defparam \Lab_UT.display.dOut_RNO_1_1_LC_9_5_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.display.dOut_RNO_1_1_LC_9_5_4 .LUT_INIT=16'b1101110011001100;
    LogicCell40 \Lab_UT.display.dOut_RNO_1_1_LC_9_5_4  (
            .in0(N__26331),
            .in1(N__26257),
            .in2(N__22882),
            .in3(N__23057),
            .lcout(\Lab_UT.display.dOutP_0_iv_i_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.display.dOut_RNO_2_3_LC_9_5_5 .C_ON=1'b0;
    defparam \Lab_UT.display.dOut_RNO_2_3_LC_9_5_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.display.dOut_RNO_2_3_LC_9_5_5 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \Lab_UT.display.dOut_RNO_2_3_LC_9_5_5  (
            .in0(_gnd_net_),
            .in1(N__26333),
            .in2(_gnd_net_),
            .in3(N__22930),
            .lcout(),
            .ltout(\Lab_UT.display.N_101_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.display.dOut_RNO_0_3_LC_9_5_6 .C_ON=1'b0;
    defparam \Lab_UT.display.dOut_RNO_0_3_LC_9_5_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.display.dOut_RNO_0_3_LC_9_5_6 .LUT_INIT=16'b1010000011101100;
    LogicCell40 \Lab_UT.display.dOut_RNO_0_3_LC_9_5_6  (
            .in0(N__22873),
            .in1(N__26540),
            .in2(N__22861),
            .in3(N__22688),
            .lcout(),
            .ltout(\Lab_UT.display.dOutP_0_iv_i_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.display.dOut_3_LC_9_5_7 .C_ON=1'b0;
    defparam \Lab_UT.display.dOut_3_LC_9_5_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.display.dOut_3_LC_9_5_7 .LUT_INIT=16'b0000000000001110;
    LogicCell40 \Lab_UT.display.dOut_3_LC_9_5_7  (
            .in0(N__23130),
            .in1(N__22858),
            .in2(N__22843),
            .in3(N__22840),
            .lcout(L3_tx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29450),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_addr_5_LC_9_6_0 .C_ON=1'b0;
    defparam \uu2.r_addr_5_LC_9_6_0 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_5_LC_9_6_0 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.r_addr_5_LC_9_6_0  (
            .in0(N__25108),
            .in1(N__25180),
            .in2(N__22792),
            .in3(N__25147),
            .lcout(\uu2.r_addrZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29442),
            .ce(),
            .sr(N__26072));
    defparam \Lab_UT.didp.Mones_alarm.q_0_LC_9_6_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mones_alarm.q_0_LC_9_6_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.Mones_alarm.q_0_LC_9_6_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Lab_UT.didp.Mones_alarm.q_0_LC_9_6_1  (
            .in0(N__22711),
            .in1(N__22760),
            .in2(_gnd_net_),
            .in3(N__29103),
            .lcout(\Lab_UT.di_AMones_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29442),
            .ce(),
            .sr(N__26072));
    defparam \Lab_UT.didp.Mones_alarm.q_1_LC_9_6_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mones_alarm.q_1_LC_9_6_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.Mones_alarm.q_1_LC_9_6_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Lab_UT.didp.Mones_alarm.q_1_LC_9_6_2  (
            .in0(N__28795),
            .in1(N__25775),
            .in2(_gnd_net_),
            .in3(N__22712),
            .lcout(\Lab_UT.di_AMones_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29442),
            .ce(),
            .sr(N__26072));
    defparam \Lab_UT.didp.Mones_alarm.q_2_LC_9_6_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mones_alarm.q_2_LC_9_6_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.Mones_alarm.q_2_LC_9_6_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Lab_UT.didp.Mones_alarm.q_2_LC_9_6_3  (
            .in0(N__22713),
            .in1(N__22734),
            .in2(_gnd_net_),
            .in3(N__28610),
            .lcout(\Lab_UT.di_AMones_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29442),
            .ce(),
            .sr(N__26072));
    defparam \Lab_UT.didp.Mones_alarm.q_3_LC_9_6_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mones_alarm.q_3_LC_9_6_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.Mones_alarm.q_3_LC_9_6_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Lab_UT.didp.Mones_alarm.q_3_LC_9_6_4  (
            .in0(N__28983),
            .in1(N__22689),
            .in2(_gnd_net_),
            .in3(N__22714),
            .lcout(\Lab_UT.di_AMones_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29442),
            .ce(),
            .sr(N__26072));
    defparam \Lab_UT.didp.Sones_alarm.q_0_LC_9_6_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.Sones_alarm.q_0_LC_9_6_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.Sones_alarm.q_0_LC_9_6_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Lab_UT.didp.Sones_alarm.q_0_LC_9_6_5  (
            .in0(N__22961),
            .in1(N__23077),
            .in2(_gnd_net_),
            .in3(N__29104),
            .lcout(\Lab_UT.di_ASones_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29442),
            .ce(),
            .sr(N__26072));
    defparam \Lab_UT.didp.Sones_alarm.q_1_LC_9_6_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.Sones_alarm.q_1_LC_9_6_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.Sones_alarm.q_1_LC_9_6_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Lab_UT.didp.Sones_alarm.q_1_LC_9_6_6  (
            .in0(N__28796),
            .in1(N__23058),
            .in2(_gnd_net_),
            .in3(N__22962),
            .lcout(\Lab_UT.di_ASones_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29442),
            .ce(),
            .sr(N__26072));
    defparam \Lab_UT.didp.Sones_alarm.q_2_LC_9_6_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.Sones_alarm.q_2_LC_9_6_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.Sones_alarm.q_2_LC_9_6_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Lab_UT.didp.Sones_alarm.q_2_LC_9_6_7  (
            .in0(N__22963),
            .in1(N__23038),
            .in2(_gnd_net_),
            .in3(N__28611),
            .lcout(\Lab_UT.di_ASones_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29442),
            .ce(),
            .sr(N__26072));
    defparam \Lab_UT.didp.Mtens_alarm.q_2_LC_9_7_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mtens_alarm.q_2_LC_9_7_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.Mtens_alarm.q_2_LC_9_7_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.didp.Mtens_alarm.q_2_LC_9_7_0  (
            .in0(N__23018),
            .in1(N__28608),
            .in2(_gnd_net_),
            .in3(N__25843),
            .lcout(\Lab_UT.di_AMtens_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29436),
            .ce(),
            .sr(N__26069));
    defparam \Lab_UT.didp.Mtens_alarm.q_3_LC_9_7_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mtens_alarm.q_3_LC_9_7_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.Mtens_alarm.q_3_LC_9_7_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Lab_UT.didp.Mtens_alarm.q_3_LC_9_7_1  (
            .in0(N__23019),
            .in1(N__25526),
            .in2(_gnd_net_),
            .in3(N__28985),
            .lcout(\Lab_UT.di_AMtens_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29436),
            .ce(),
            .sr(N__26069));
    defparam \Lab_UT.didp.Stens_alarm.q_2_LC_9_7_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.Stens_alarm.q_2_LC_9_7_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.Stens_alarm.q_2_LC_9_7_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \Lab_UT.didp.Stens_alarm.q_2_LC_9_7_2  (
            .in0(N__25629),
            .in1(N__28609),
            .in2(_gnd_net_),
            .in3(N__22908),
            .lcout(\Lab_UT.di_AStens_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29436),
            .ce(),
            .sr(N__26069));
    defparam \Lab_UT.didp.Stens_alarm.q_3_LC_9_7_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.Stens_alarm.q_3_LC_9_7_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.Stens_alarm.q_3_LC_9_7_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Lab_UT.didp.Stens_alarm.q_3_LC_9_7_3  (
            .in0(N__22909),
            .in1(N__22983),
            .in2(_gnd_net_),
            .in3(N__28986),
            .lcout(\Lab_UT.di_AStens_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29436),
            .ce(),
            .sr(N__26069));
    defparam \Lab_UT.didp.Sones_alarm.q_3_LC_9_7_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.Sones_alarm.q_3_LC_9_7_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.Sones_alarm.q_3_LC_9_7_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Lab_UT.didp.Sones_alarm.q_3_LC_9_7_4  (
            .in0(N__28984),
            .in1(N__22953),
            .in2(_gnd_net_),
            .in3(N__22929),
            .lcout(\Lab_UT.di_ASones_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29436),
            .ce(),
            .sr(N__26069));
    defparam \Lab_UT.didp.Stens_alarm.q_0_LC_9_7_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.Stens_alarm.q_0_LC_9_7_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.Stens_alarm.q_0_LC_9_7_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Lab_UT.didp.Stens_alarm.q_0_LC_9_7_5  (
            .in0(N__22906),
            .in1(N__25728),
            .in2(_gnd_net_),
            .in3(N__29105),
            .lcout(\Lab_UT.di_AStens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29436),
            .ce(),
            .sr(N__26069));
    defparam \Lab_UT.didp.Stens_alarm.q_1_LC_9_7_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.Stens_alarm.q_1_LC_9_7_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.Stens_alarm.q_1_LC_9_7_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Lab_UT.didp.Stens_alarm.q_1_LC_9_7_6  (
            .in0(N__28816),
            .in1(N__25802),
            .in2(_gnd_net_),
            .in3(N__22907),
            .lcout(\Lab_UT.di_AStens_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29436),
            .ce(),
            .sr(N__26069));
    defparam \Lab_UT.uu0.sec_clk_LC_9_7_7 .C_ON=1'b0;
    defparam \Lab_UT.uu0.sec_clk_LC_9_7_7 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.uu0.sec_clk_LC_9_7_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \Lab_UT.uu0.sec_clk_LC_9_7_7  (
            .in0(N__23246),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23157),
            .lcout(\Lab_UT.halfPulse ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29436),
            .ce(),
            .sr(N__26069));
    defparam \Lab_UT.didp.Stens_subtractor.q_7_i_o2_2_LC_9_8_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.Stens_subtractor.q_7_i_o2_2_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Stens_subtractor.q_7_i_o2_2_LC_9_8_0 .LUT_INIT=16'b0101110101111111;
    LogicCell40 \Lab_UT.didp.Stens_subtractor.q_7_i_o2_2_LC_9_8_0  (
            .in0(N__28180),
            .in1(N__29959),
            .in2(N__23112),
            .in3(N__23091),
            .lcout(\Lab_UT.didp.Stens_subtractor.N_86 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.displayAlarm_1_LC_9_8_1 .C_ON=1'b0;
    defparam \Lab_UT.displayAlarm_1_LC_9_8_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.displayAlarm_1_LC_9_8_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.displayAlarm_1_LC_9_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29540),
            .lcout(\Lab_UT.displayAlarmZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29427),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.dicLdStens_RNIQVHE3_LC_9_8_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.dicLdStens_RNIQVHE3_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.dicLdStens_RNIQVHE3_LC_9_8_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Lab_UT.dictrl.dicLdStens_RNIQVHE3_LC_9_8_2  (
            .in0(N__23105),
            .in1(N__29958),
            .in2(_gnd_net_),
            .in3(N__23090),
            .lcout(\Lab_UT.ld_enable_Stens ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Stens_subtractor.q_RNI8PD76_1_LC_9_8_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.Stens_subtractor.q_RNI8PD76_1_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Stens_subtractor.q_RNI8PD76_1_LC_9_8_3 .LUT_INIT=16'b1110111000010001;
    LogicCell40 \Lab_UT.didp.Stens_subtractor.q_RNI8PD76_1_LC_9_8_3  (
            .in0(N__26620),
            .in1(N__29683),
            .in2(_gnd_net_),
            .in3(N__27873),
            .lcout(\Lab_UT.didp.Stens_subtractor.q_RNI8PD76Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Stens_subtractor.q_RNIBBF11_2_LC_9_8_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.Stens_subtractor.q_RNIBBF11_2_LC_9_8_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Stens_subtractor.q_RNIBBF11_2_LC_9_8_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \Lab_UT.didp.Stens_subtractor.q_RNIBBF11_2_LC_9_8_4  (
            .in0(N__26233),
            .in1(N__29761),
            .in2(_gnd_net_),
            .in3(N__27161),
            .lcout(\Lab_UT.didp.q_RNIBBF11_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Stens_subtractor.q_RNO_0_3_LC_9_8_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.Stens_subtractor.q_RNO_0_3_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Stens_subtractor.q_RNO_0_3_LC_9_8_5 .LUT_INIT=16'b0110110011001001;
    LogicCell40 \Lab_UT.didp.Stens_subtractor.q_RNO_0_3_LC_9_8_5  (
            .in0(N__26623),
            .in1(N__27118),
            .in2(N__26602),
            .in3(N__27159),
            .lcout(\Lab_UT.didp.Stens_subtractor.q_RNO_0_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Stens_subtractor.q_RNO_0_2_LC_9_8_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.Stens_subtractor.q_RNO_0_2_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Stens_subtractor.q_RNO_0_2_LC_9_8_6 .LUT_INIT=16'b1111111000000001;
    LogicCell40 \Lab_UT.didp.Stens_subtractor.q_RNO_0_2_LC_9_8_6  (
            .in0(N__29685),
            .in1(N__26622),
            .in2(N__27877),
            .in3(N__27160),
            .lcout(\Lab_UT.didp.Stens_subtractor.q_RNO_0_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Stens_subtractor.q_RNO_0_0_LC_9_8_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.Stens_subtractor.q_RNO_0_0_LC_9_8_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Stens_subtractor.q_RNO_0_0_LC_9_8_7 .LUT_INIT=16'b1001100110011001;
    LogicCell40 \Lab_UT.didp.Stens_subtractor.q_RNO_0_0_LC_9_8_7  (
            .in0(N__26621),
            .in1(N__29684),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.didp.Stens_subtractor.un1_q_axb0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Stens_subtractor.q_0_LC_9_9_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.Stens_subtractor.q_0_LC_9_9_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.Stens_subtractor.q_0_LC_9_9_0 .LUT_INIT=16'b1111110101110101;
    LogicCell40 \Lab_UT.didp.Stens_subtractor.q_0_LC_9_9_0  (
            .in0(N__26969),
            .in1(N__23549),
            .in2(N__29106),
            .in3(N__23563),
            .lcout(\Lab_UT.didp.di_Stens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29417),
            .ce(),
            .sr(N__28448));
    defparam \Lab_UT.didp.Stens_subtractor.q_3_LC_9_9_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.Stens_subtractor.q_3_LC_9_9_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.Stens_subtractor.q_3_LC_9_9_1 .LUT_INIT=16'b1101100000000000;
    LogicCell40 \Lab_UT.didp.Stens_subtractor.q_3_LC_9_9_1  (
            .in0(N__23551),
            .in1(N__23557),
            .in2(N__28995),
            .in3(N__26971),
            .lcout(\Lab_UT.didp.di_Stens_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29417),
            .ce(),
            .sr(N__28448));
    defparam \Lab_UT.didp.Stens_subtractor.q_2_LC_9_9_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.Stens_subtractor.q_2_LC_9_9_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.Stens_subtractor.q_2_LC_9_9_2 .LUT_INIT=16'b1111110101110101;
    LogicCell40 \Lab_UT.didp.Stens_subtractor.q_2_LC_9_9_2  (
            .in0(N__26970),
            .in1(N__23550),
            .in2(N__28612),
            .in3(N__23539),
            .lcout(\Lab_UT.didp.di_Stens_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29417),
            .ce(),
            .sr(N__28448));
    defparam \Lab_UT.didp.Stens_subtractor.q_RNIDDF11_3_LC_9_9_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.Stens_subtractor.q_RNIDDF11_3_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Stens_subtractor.q_RNIDDF11_3_LC_9_9_3 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \Lab_UT.didp.Stens_subtractor.q_RNIDDF11_3_LC_9_9_3  (
            .in0(N__27119),
            .in1(_gnd_net_),
            .in2(N__29779),
            .in3(N__26197),
            .lcout(),
            .ltout(\Lab_UT.didp.q_RNIDDF11_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.curr_LED_RNIRNM52_1_LC_9_9_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.curr_LED_RNIRNM52_1_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.curr_LED_RNIRNM52_1_LC_9_9_4 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \Lab_UT.didp.curr_LED_RNIRNM52_1_LC_9_9_4  (
            .in0(N__29630),
            .in1(_gnd_net_),
            .in2(N__23533),
            .in3(N__23518),
            .lcout(led_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Mones_subtractor.q_RNI1TVP_3_LC_9_9_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mones_subtractor.q_RNI1TVP_3_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Mones_subtractor.q_RNI1TVP_3_LC_9_9_5 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \Lab_UT.didp.Mones_subtractor.q_RNI1TVP_3_LC_9_9_5  (
            .in0(N__26832),
            .in1(_gnd_net_),
            .in2(N__29778),
            .in3(N__28252),
            .lcout(\Lab_UT.didp.q_RNI1TVP_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.curr_LED_RNINJM52_1_LC_9_9_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.curr_LED_RNINJM52_1_LC_9_9_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.curr_LED_RNINJM52_1_LC_9_9_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \Lab_UT.didp.curr_LED_RNINJM52_1_LC_9_9_7  (
            .in0(N__23512),
            .in1(N__23506),
            .in2(_gnd_net_),
            .in3(N__29629),
            .lcout(led_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.r_dicRun_LC_9_10_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.r_dicRun_LC_9_10_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.r_dicRun_LC_9_10_0 .LUT_INIT=16'b0100010000000101;
    LogicCell40 \Lab_UT.dictrl.r_dicRun_LC_9_10_0  (
            .in0(N__23482),
            .in1(N__26667),
            .in2(N__24742),
            .in3(N__23456),
            .lcout(\Lab_UT.ld_enable_dicRun ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29410),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_al_0_LC_9_10_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_al_0_LC_9_10_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.nextState_al_0_LC_9_10_1 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \Lab_UT.dictrl.nextState_al_0_LC_9_10_1  (
            .in0(N__23572),
            .in1(N__23605),
            .in2(N__24121),
            .in3(N__26156),
            .lcout(\Lab_UT.dictrl.nextState_al_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29410),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.r_dicAlarmArmed_LC_9_10_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.r_dicAlarmArmed_LC_9_10_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.r_dicAlarmArmed_LC_9_10_2 .LUT_INIT=16'b0010000000110011;
    LogicCell40 \Lab_UT.dictrl.r_dicAlarmArmed_LC_9_10_2  (
            .in0(N__29576),
            .in1(N__29126),
            .in2(N__27395),
            .in3(N__24058),
            .lcout(\Lab_UT.alarm_armed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29410),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.r_dicAlarmTrig_LC_9_10_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.r_dicAlarmTrig_LC_9_10_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.r_dicAlarmTrig_LC_9_10_3 .LUT_INIT=16'b0000111000000010;
    LogicCell40 \Lab_UT.dictrl.r_dicAlarmTrig_LC_9_10_3  (
            .in0(N__24057),
            .in1(N__29577),
            .in2(N__29130),
            .in3(N__23645),
            .lcout(\Lab_UT.dictrl.r_dicAlarmTrigZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29410),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.displayAlarm_5_LC_9_10_5 .C_ON=1'b0;
    defparam \Lab_UT.displayAlarm_5_LC_9_10_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.displayAlarm_5_LC_9_10_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Lab_UT.displayAlarm_5_LC_9_10_5  (
            .in0(_gnd_net_),
            .in1(N__29539),
            .in2(_gnd_net_),
            .in3(N__27388),
            .lcout(\Lab_UT.displayAlarmZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29410),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_al_RNIHVQHE_0_LC_9_10_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_al_RNIHVQHE_0_LC_9_10_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_al_RNIHVQHE_0_LC_9_10_6 .LUT_INIT=16'b1111010110110001;
    LogicCell40 \Lab_UT.dictrl.nextState_al_RNIHVQHE_0_LC_9_10_6  (
            .in0(N__29575),
            .in1(N__24084),
            .in2(N__24120),
            .in3(N__24133),
            .lcout(\Lab_UT.dictrl.nextState_al_1 ),
            .ltout(\Lab_UT.dictrl.nextState_al_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_al_ret_LC_9_10_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_al_ret_LC_9_10_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.currState_al_ret_LC_9_10_7 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \Lab_UT.dictrl.currState_al_ret_LC_9_10_7  (
            .in0(N__23571),
            .in1(_gnd_net_),
            .in2(N__23599),
            .in3(N__26157),
            .lcout(\Lab_UT.dictrl.un1_nextState_al24_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29410),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_al_0_0_LC_9_11_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_al_0_0_LC_9_11_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.currState_al_0_0_LC_9_11_0 .LUT_INIT=16'b1101000111000000;
    LogicCell40 \Lab_UT.dictrl.currState_al_0_0_LC_9_11_0  (
            .in0(N__24055),
            .in1(N__29573),
            .in2(N__24127),
            .in3(N__23581),
            .lcout(\Lab_UT.dictrl.currState_alZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29403),
            .ce(),
            .sr(N__26073));
    defparam \Lab_UT.dictrl.currState_al_0_RNIRBNK8_0_LC_9_11_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_al_0_RNIRBNK8_0_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_al_0_RNIRBNK8_0_LC_9_11_1 .LUT_INIT=16'b0000101110111011;
    LogicCell40 \Lab_UT.dictrl.currState_al_0_RNIRBNK8_0_LC_9_11_1  (
            .in0(N__24496),
            .in1(N__24052),
            .in2(N__24073),
            .in3(N__27355),
            .lcout(\Lab_UT.dictrl.nextState_al_1_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_0_ret_15_RNILDPC8_LC_9_11_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_15_RNILDPC8_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_0_ret_15_RNILDPC8_LC_9_11_2 .LUT_INIT=16'b0011000101000100;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_15_RNILDPC8_LC_9_11_2  (
            .in0(N__27354),
            .in1(N__24068),
            .in2(N__23596),
            .in3(N__24495),
            .lcout(\Lab_UT.dictrl.nextState_al_latmux_1 ),
            .ltout(\Lab_UT.dictrl.nextState_al_latmux_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.nextState_al_RNISS2D9_0_LC_9_11_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.nextState_al_RNISS2D9_0_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.nextState_al_RNISS2D9_0_LC_9_11_3 .LUT_INIT=16'b1000100011011000;
    LogicCell40 \Lab_UT.dictrl.nextState_al_RNISS2D9_0_LC_9_11_3  (
            .in0(N__29572),
            .in1(N__24122),
            .in2(N__23575),
            .in3(N__24054),
            .lcout(\Lab_UT.dictrl.nextState_alZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_al_0_RNI5PG55_1_LC_9_11_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_al_0_RNI5PG55_1_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_al_0_RNI5PG55_1_LC_9_11_5 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \Lab_UT.dictrl.currState_al_0_RNI5PG55_1_LC_9_11_5  (
            .in0(N__24056),
            .in1(N__27353),
            .in2(_gnd_net_),
            .in3(N__24178),
            .lcout(\Lab_UT.dictrl.N_186 ),
            .ltout(\Lab_UT.dictrl.N_186_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_al_0_1_LC_9_11_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_al_0_1_LC_9_11_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.currState_al_0_1_LC_9_11_6 .LUT_INIT=16'b1011100010111011;
    LogicCell40 \Lab_UT.dictrl.currState_al_0_1_LC_9_11_6  (
            .in0(N__24126),
            .in1(N__29574),
            .in2(N__24088),
            .in3(N__24085),
            .lcout(\Lab_UT.dictrl.currState_alZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29403),
            .ce(),
            .sr(N__26073));
    defparam \Lab_UT.dictrl.currState_al_0_RNIB8DH_0_LC_9_11_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_al_0_RNIB8DH_0_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_al_0_RNIB8DH_0_LC_9_11_7 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \Lab_UT.dictrl.currState_al_0_RNIB8DH_0_LC_9_11_7  (
            .in0(N__24072),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24053),
            .lcout(\Lab_UT.dictrl.nextState_al22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_0_ret_0_RNIHG3F_LC_9_12_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_0_RNIHG3F_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_0_ret_0_RNIHG3F_LC_9_12_0 .LUT_INIT=16'b0010111011101110;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_0_RNIHG3F_LC_9_12_0  (
            .in0(N__23855),
            .in1(N__23777),
            .in2(N__24028),
            .in3(N__24013),
            .lcout(),
            .ltout(\Lab_UT.dictrl.un1_currState_8_u_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_ret_7_RNI03VH1_LC_9_12_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_ret_7_RNI03VH1_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_ret_7_RNI03VH1_LC_9_12_1 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \Lab_UT.dictrl.currState_ret_7_RNI03VH1_LC_9_12_1  (
            .in0(N__24886),
            .in1(N__24514),
            .in2(N__23923),
            .in3(N__25023),
            .lcout(\Lab_UT.dictrl.currState_ret_7_RNI03VHZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_ret_7_RNI2HHP_LC_9_12_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_ret_7_RNI2HHP_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_ret_7_RNI2HHP_LC_9_12_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.dictrl.currState_ret_7_RNI2HHP_LC_9_12_2  (
            .in0(_gnd_net_),
            .in1(N__24512),
            .in2(_gnd_net_),
            .in3(N__24885),
            .lcout(\Lab_UT.dictrl.un1_currState_inv_1 ),
            .ltout(\Lab_UT.dictrl.un1_currState_inv_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_0_ret_1_RNIPH7F1_LC_9_12_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_1_RNIPH7F1_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_0_ret_1_RNIPH7F1_LC_9_12_3 .LUT_INIT=16'b1111000001100110;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_1_RNIPH7F1_LC_9_12_3  (
            .in0(N__23775),
            .in1(N__23856),
            .in2(N__23902),
            .in3(N__25021),
            .lcout(\Lab_UT.dictrl.currState_0_ret_1_RNIPH7FZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_0_ret_5_RNI9PAE_LC_9_12_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_5_RNI9PAE_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_0_ret_5_RNI9PAE_LC_9_12_4 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_5_RNI9PAE_LC_9_12_4  (
            .in0(N__23869),
            .in1(N__23854),
            .in2(_gnd_net_),
            .in3(N__23776),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_201_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_2_RNIOB6H1_2_LC_9_12_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_2_RNIOB6H1_2_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_2_RNIOB6H1_2_LC_9_12_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \Lab_UT.dictrl.currState_2_RNIOB6H1_2_LC_9_12_5  (
            .in0(_gnd_net_),
            .in1(N__23685),
            .in2(N__23674),
            .in3(N__25022),
            .lcout(\Lab_UT.dictrl.currState_2_RNIOB6H1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.r_dicRun_RNO_0_LC_9_12_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.r_dicRun_RNO_0_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.r_dicRun_RNO_0_LC_9_12_6 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \Lab_UT.dictrl.r_dicRun_RNO_0_LC_9_12_6  (
            .in0(N__25024),
            .in1(N__24513),
            .in2(_gnd_net_),
            .in3(N__24887),
            .lcout(\Lab_UT.dictrl.r_dicRun_r_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_ret_7_LC_9_12_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_ret_7_LC_9_12_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.currState_ret_7_LC_9_12_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Lab_UT.dictrl.currState_ret_7_LC_9_12_7  (
            .in0(_gnd_net_),
            .in1(N__24725),
            .in2(_gnd_net_),
            .in3(N__24706),
            .lcout(\Lab_UT.dictrl.r_dicLdMtens15_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29397),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.decoder.de_atSign_4_LC_9_13_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.decoder.de_atSign_4_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.decoder.de_atSign_4_LC_9_13_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \Lab_UT.dictrl.decoder.de_atSign_4_LC_9_13_0  (
            .in0(N__24446),
            .in1(N__29062),
            .in2(N__24322),
            .in3(N__28539),
            .lcout(),
            .ltout(\Lab_UT.dictrl.decoder.de_atSignZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.decoder.de_atSign_LC_9_13_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.decoder.de_atSign_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.decoder.de_atSign_LC_9_13_1 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \Lab_UT.dictrl.decoder.de_atSign_LC_9_13_1  (
            .in0(_gnd_net_),
            .in1(N__25225),
            .in2(N__24499),
            .in3(N__27794),
            .lcout(\Lab_UT.dictrl.de_atSign ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.decoder.de_littleA_2_LC_9_13_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.decoder.de_littleA_2_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.decoder.de_littleA_2_LC_9_13_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \Lab_UT.dictrl.decoder.de_littleA_2_LC_9_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24321),
            .in3(N__24444),
            .lcout(\Lab_UT.dictrl.de_littleA_2 ),
            .ltout(\Lab_UT.dictrl.de_littleA_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.decoder.de_littleL_LC_9_13_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.decoder.de_littleL_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.decoder.de_littleL_LC_9_13_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.decoder.de_littleL_LC_9_13_3  (
            .in0(N__25490),
            .in1(N__24347),
            .in2(N__24484),
            .in3(N__27793),
            .lcout(\Lab_UT.dictrl.de_littleL ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.decoder.g0_4_2_LC_9_13_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.decoder.g0_4_2_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.decoder.g0_4_2_LC_9_13_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.decoder.g0_4_2_LC_9_13_4  (
            .in0(N__24445),
            .in1(N__24340),
            .in2(N__24320),
            .in3(N__25489),
            .lcout(\Lab_UT.dictrl.g0_4_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.decoder.de_littleN_1_LC_9_13_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.decoder.de_littleN_1_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.decoder.de_littleN_1_LC_9_13_5 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \Lab_UT.dictrl.decoder.de_littleN_1_LC_9_13_5  (
            .in0(N__29064),
            .in1(N__28756),
            .in2(N__24206),
            .in3(N__25315),
            .lcout(),
            .ltout(\Lab_UT.dictrl.decoder.de_littleNZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.decoder.de_littleN_LC_9_13_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.decoder.de_littleN_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.decoder.de_littleN_LC_9_13_6 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \Lab_UT.dictrl.decoder.de_littleN_LC_9_13_6  (
            .in0(N__27795),
            .in1(N__25402),
            .in2(N__25495),
            .in3(N__25491),
            .lcout(\Lab_UT.n_rdy ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.escKey_3_LC_9_13_7 .C_ON=1'b0;
    defparam \resetGen.escKey_3_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \resetGen.escKey_3_LC_9_13_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \resetGen.escKey_3_LC_9_13_7  (
            .in0(N__29063),
            .in1(N__28755),
            .in2(N__28994),
            .in3(N__25314),
            .lcout(\resetGen.escKeyZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_1_LC_9_14_3 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_1_LC_9_14_3 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_1_LC_9_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_1_LC_9_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28563),
            .lcout(bu_rx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29387),
            .ce(N__25427),
            .sr(N__26103));
    defparam \buart.Z_rx.shifter_2_LC_9_14_6 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_2_LC_9_14_6 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_2_LC_9_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_2_LC_9_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28905),
            .lcout(bu_rx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29387),
            .ce(N__25427),
            .sr(N__26103));
    defparam \Lab_UT.dictrl.decoder.de_atSign_5_LC_9_15_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.decoder.de_atSign_5_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.decoder.de_atSign_5_LC_9_15_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Lab_UT.dictrl.decoder.de_atSign_5_LC_9_15_1  (
            .in0(N__28754),
            .in1(N__25376),
            .in2(N__28943),
            .in3(N__25313),
            .lcout(\Lab_UT.dictrl.decoder.de_atSignZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.uu0.l_precount_0_LC_11_2_5 .C_ON=1'b0;
    defparam \Lab_UT.uu0.l_precount_0_LC_11_2_5 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.uu0.l_precount_0_LC_11_2_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Lab_UT.uu0.l_precount_0_LC_11_2_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25199),
            .lcout(\Lab_UT.uu0.l_precountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29477),
            .ce(),
            .sr(N__26106));
    defparam \uu2.r_addr_4_LC_11_3_6 .C_ON=1'b0;
    defparam \uu2.r_addr_4_LC_11_3_6 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_4_LC_11_3_6 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \uu2.r_addr_4_LC_11_3_6  (
            .in0(N__25088),
            .in1(N__25179),
            .in2(_gnd_net_),
            .in3(N__25146),
            .lcout(\uu2.r_addrZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29473),
            .ce(),
            .sr(N__26075));
    defparam \Lab_UT.displayAlarm_0_LC_11_4_0 .C_ON=1'b0;
    defparam \Lab_UT.displayAlarm_0_LC_11_4_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.displayAlarm_0_LC_11_4_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.displayAlarm_0_LC_11_4_0  (
            .in0(_gnd_net_),
            .in1(N__29548),
            .in2(_gnd_net_),
            .in3(N__27414),
            .lcout(\Lab_UT.displayAlarmZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29466),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.display.dOut_RNO_2_0_LC_11_4_1 .C_ON=1'b0;
    defparam \Lab_UT.display.dOut_RNO_2_0_LC_11_4_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.display.dOut_RNO_2_0_LC_11_4_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Lab_UT.display.dOut_RNO_2_0_LC_11_4_1  (
            .in0(_gnd_net_),
            .in1(N__25867),
            .in2(_gnd_net_),
            .in3(N__25069),
            .lcout(\Lab_UT.display.N_130 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.display.dOut_RNO_0_0_LC_11_4_2 .C_ON=1'b0;
    defparam \Lab_UT.display.dOut_RNO_0_0_LC_11_4_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.display.dOut_RNO_0_0_LC_11_4_2 .LUT_INIT=16'b0000110010101110;
    LogicCell40 \Lab_UT.display.dOut_RNO_0_0_LC_11_4_2  (
            .in0(N__25659),
            .in1(N__25875),
            .in2(N__25741),
            .in3(N__25732),
            .lcout(),
            .ltout(\Lab_UT.display.dOutP_0_iv_i_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.display.dOut_0_LC_11_4_3 .C_ON=1'b0;
    defparam \Lab_UT.display.dOut_0_LC_11_4_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.display.dOut_0_LC_11_4_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Lab_UT.display.dOut_0_LC_11_4_3  (
            .in0(N__26439),
            .in1(N__25708),
            .in2(N__25702),
            .in3(N__25699),
            .lcout(L3_tx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29466),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.displayAlarm_2_LC_11_4_4 .C_ON=1'b0;
    defparam \Lab_UT.displayAlarm_2_LC_11_4_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.displayAlarm_2_LC_11_4_4 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \Lab_UT.displayAlarm_2_LC_11_4_4  (
            .in0(_gnd_net_),
            .in1(N__29547),
            .in2(_gnd_net_),
            .in3(N__27415),
            .lcout(\Lab_UT.displayAlarmZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29466),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.display.dOut_RNO_0_2_LC_11_4_5 .C_ON=1'b0;
    defparam \Lab_UT.display.dOut_RNO_0_2_LC_11_4_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.display.dOut_RNO_0_2_LC_11_4_5 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \Lab_UT.display.dOut_RNO_0_2_LC_11_4_5  (
            .in0(N__25876),
            .in1(N__25660),
            .in2(N__25645),
            .in3(N__25633),
            .lcout(),
            .ltout(\Lab_UT.display.dOutP_0_iv_i_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.display.dOut_2_LC_11_4_6 .C_ON=1'b0;
    defparam \Lab_UT.display.dOut_2_LC_11_4_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.display.dOut_2_LC_11_4_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Lab_UT.display.dOut_2_LC_11_4_6  (
            .in0(N__25816),
            .in1(N__26440),
            .in2(N__25609),
            .in3(N__25606),
            .lcout(L3_tx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29466),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.display.cnt_RNIFA8M_2_LC_11_4_7 .C_ON=1'b0;
    defparam \Lab_UT.display.cnt_RNIFA8M_2_LC_11_4_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.display.cnt_RNIFA8M_2_LC_11_4_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Lab_UT.display.cnt_RNIFA8M_2_LC_11_4_7  (
            .in0(N__26406),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26486),
            .lcout(\Lab_UT.display.un42_dOutP_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.display.cnt_RNI1STE1_1_LC_11_5_0 .C_ON=1'b0;
    defparam \Lab_UT.display.cnt_RNI1STE1_1_LC_11_5_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.display.cnt_RNI1STE1_1_LC_11_5_0 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \Lab_UT.display.cnt_RNI1STE1_1_LC_11_5_0  (
            .in0(N__25865),
            .in1(N__26496),
            .in2(_gnd_net_),
            .in3(N__26732),
            .lcout(\Lab_UT.display.cnt_RNI1STE1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.display.cnt_RNIE98M_2_LC_11_5_1 .C_ON=1'b0;
    defparam \Lab_UT.display.cnt_RNIE98M_2_LC_11_5_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.display.cnt_RNIE98M_2_LC_11_5_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Lab_UT.display.cnt_RNIE98M_2_LC_11_5_1  (
            .in0(_gnd_net_),
            .in1(N__26401),
            .in2(_gnd_net_),
            .in3(N__26297),
            .lcout(\Lab_UT.display.N_151 ),
            .ltout(\Lab_UT.display.N_151_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.display.dOut_RNO_3_3_LC_11_5_2 .C_ON=1'b0;
    defparam \Lab_UT.display.dOut_RNO_3_3_LC_11_5_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.display.dOut_RNO_3_3_LC_11_5_2 .LUT_INIT=16'b0001000001010000;
    LogicCell40 \Lab_UT.display.dOut_RNO_3_3_LC_11_5_2  (
            .in0(N__26501),
            .in1(N__26731),
            .in2(N__25537),
            .in3(N__25534),
            .lcout(\Lab_UT.display.N_124 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.display.cnt_0_LC_11_5_3 .C_ON=1'b0;
    defparam \Lab_UT.display.cnt_0_LC_11_5_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.display.cnt_0_LC_11_5_3 .LUT_INIT=16'b0000000011111110;
    LogicCell40 \Lab_UT.display.cnt_0_LC_11_5_3  (
            .in0(N__26733),
            .in1(N__26402),
            .in2(N__26510),
            .in3(N__26300),
            .lcout(\Lab_UT.display.cntZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29458),
            .ce(),
            .sr(N__26074));
    defparam \Lab_UT.display.cnt_2_LC_11_5_4 .C_ON=1'b0;
    defparam \Lab_UT.display.cnt_2_LC_11_5_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.display.cnt_2_LC_11_5_4 .LUT_INIT=16'b0101101011110000;
    LogicCell40 \Lab_UT.display.cnt_2_LC_11_5_4  (
            .in0(N__26299),
            .in1(_gnd_net_),
            .in2(N__26417),
            .in3(N__26500),
            .lcout(\Lab_UT.display.cntZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29458),
            .ce(),
            .sr(N__26074));
    defparam \Lab_UT.display.cnt_1_LC_11_5_5 .C_ON=1'b0;
    defparam \Lab_UT.display.cnt_1_LC_11_5_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.display.cnt_1_LC_11_5_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Lab_UT.display.cnt_1_LC_11_5_5  (
            .in0(_gnd_net_),
            .in1(N__26502),
            .in2(_gnd_net_),
            .in3(N__26301),
            .lcout(\Lab_UT.display.cntZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29458),
            .ce(),
            .sr(N__26074));
    defparam \Lab_UT.display.cnt_RNID88M_1_LC_11_5_6 .C_ON=1'b0;
    defparam \Lab_UT.display.cnt_RNID88M_1_LC_11_5_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.display.cnt_RNID88M_1_LC_11_5_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Lab_UT.display.cnt_RNID88M_1_LC_11_5_6  (
            .in0(N__26298),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26495),
            .lcout(\Lab_UT.display.N_106 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.display.dOut_RNO_2_2_LC_11_5_7 .C_ON=1'b0;
    defparam \Lab_UT.display.dOut_RNO_2_2_LC_11_5_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.display.dOut_RNO_2_2_LC_11_5_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Lab_UT.display.dOut_RNO_2_2_LC_11_5_7  (
            .in0(_gnd_net_),
            .in1(N__25866),
            .in2(_gnd_net_),
            .in3(N__25851),
            .lcout(\Lab_UT.display.N_115 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Stens_subtractor.q_1_LC_11_6_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.Stens_subtractor.q_1_LC_11_6_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.Stens_subtractor.q_1_LC_11_6_0 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \Lab_UT.didp.Stens_subtractor.q_1_LC_11_6_0  (
            .in0(N__26590),
            .in1(N__26551),
            .in2(N__26960),
            .in3(N__26569),
            .lcout(\Lab_UT.didp.di_Stens_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29451),
            .ce(),
            .sr(N__28419));
    defparam \Lab_UT.didp.Mones_subtractor.q_RNI775L5_3_LC_11_6_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mones_subtractor.q_RNI775L5_3_LC_11_6_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Mones_subtractor.q_RNI775L5_3_LC_11_6_2 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \Lab_UT.didp.Mones_subtractor.q_RNI775L5_3_LC_11_6_2  (
            .in0(N__26950),
            .in1(N__28024),
            .in2(_gnd_net_),
            .in3(N__27052),
            .lcout(\Lab_UT.didp.Mones_subtractor.N_80 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.display.dOut_RNO_2_1_LC_11_6_3 .C_ON=1'b0;
    defparam \Lab_UT.display.dOut_RNO_2_1_LC_11_6_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.display.dOut_RNO_2_1_LC_11_6_3 .LUT_INIT=16'b0100010100000000;
    LogicCell40 \Lab_UT.display.dOut_RNO_2_1_LC_11_6_3  (
            .in0(N__26407),
            .in1(N__25810),
            .in2(N__26334),
            .in3(N__26491),
            .lcout(),
            .ltout(\Lab_UT.display.N_108_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.display.dOut_RNO_0_1_LC_11_6_4 .C_ON=1'b0;
    defparam \Lab_UT.display.dOut_RNO_0_1_LC_11_6_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.display.dOut_RNO_0_1_LC_11_6_4 .LUT_INIT=16'b1111001011110000;
    LogicCell40 \Lab_UT.display.dOut_RNO_0_1_LC_11_6_4  (
            .in0(N__26526),
            .in1(N__26409),
            .in2(N__25783),
            .in3(N__25779),
            .lcout(\Lab_UT.display.dOutP_0_iv_i_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.display.cnt_RNID88M_0_1_LC_11_6_5 .C_ON=1'b0;
    defparam \Lab_UT.display.cnt_RNID88M_0_1_LC_11_6_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.display.cnt_RNID88M_0_1_LC_11_6_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.display.cnt_RNID88M_0_1_LC_11_6_5  (
            .in0(_gnd_net_),
            .in1(N__26490),
            .in2(_gnd_net_),
            .in3(N__26292),
            .lcout(\Lab_UT.display.N_152 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.display.cnt_RNI1STE1_2_LC_11_6_6 .C_ON=1'b0;
    defparam \Lab_UT.display.cnt_RNI1STE1_2_LC_11_6_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.display.cnt_RNI1STE1_2_LC_11_6_6 .LUT_INIT=16'b0011000000001101;
    LogicCell40 \Lab_UT.display.cnt_RNI1STE1_2_LC_11_6_6  (
            .in0(N__26730),
            .in1(N__26503),
            .in2(N__26317),
            .in3(N__26410),
            .lcout(\Lab_UT.display.N_92 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.display.dOut_RNO_3_1_LC_11_6_7 .C_ON=1'b0;
    defparam \Lab_UT.display.dOut_RNO_3_1_LC_11_6_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.display.dOut_RNO_3_1_LC_11_6_7 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \Lab_UT.display.dOut_RNO_3_1_LC_11_6_7  (
            .in0(N__26408),
            .in1(N__26729),
            .in2(N__26365),
            .in3(N__26293),
            .lcout(\Lab_UT.display.N_112 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Sones_subtractor.q_RNO_0_3_LC_11_7_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.Sones_subtractor.q_RNO_0_3_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Sones_subtractor.q_RNO_0_3_LC_11_7_0 .LUT_INIT=16'b0111100011100001;
    LogicCell40 \Lab_UT.didp.Sones_subtractor.q_RNO_0_3_LC_11_7_0  (
            .in0(N__28197),
            .in1(N__26225),
            .in2(N__26193),
            .in3(N__28030),
            .lcout(),
            .ltout(\Lab_UT.didp.Sones_subtractor.q_RNO_0Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Sones_subtractor.q_3_LC_11_7_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.Sones_subtractor.q_3_LC_11_7_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.Sones_subtractor.q_3_LC_11_7_1 .LUT_INIT=16'b1111011111010101;
    LogicCell40 \Lab_UT.didp.Sones_subtractor.q_3_LC_11_7_1  (
            .in0(N__28171),
            .in1(N__28126),
            .in2(N__26245),
            .in3(N__28996),
            .lcout(\Lab_UT.didp.di_Sones_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29443),
            .ce(),
            .sr(N__28436));
    defparam \Lab_UT.didp.Sones_subtractor.q_2_LC_11_7_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.Sones_subtractor.q_2_LC_11_7_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.Sones_subtractor.q_2_LC_11_7_2 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \Lab_UT.didp.Sones_subtractor.q_2_LC_11_7_2  (
            .in0(N__28615),
            .in1(N__28125),
            .in2(N__26242),
            .in3(N__28172),
            .lcout(\Lab_UT.didp.di_Sones_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29443),
            .ce(),
            .sr(N__28436));
    defparam \Lab_UT.didp.Sones_subtractor.q_RNO_0_2_LC_11_7_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.Sones_subtractor.q_RNO_0_2_LC_11_7_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Sones_subtractor.q_RNO_0_2_LC_11_7_3 .LUT_INIT=16'b1100110011001001;
    LogicCell40 \Lab_UT.didp.Sones_subtractor.q_RNO_0_2_LC_11_7_3  (
            .in0(N__29813),
            .in1(N__26224),
            .in2(N__28102),
            .in3(N__28196),
            .lcout(\Lab_UT.didp.Sones_subtractor.q_RNO_0_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Sones_subtractor.q_RNIIFEO1_3_LC_11_7_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.Sones_subtractor.q_RNIIFEO1_3_LC_11_7_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Sones_subtractor.q_RNIIFEO1_3_LC_11_7_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Lab_UT.didp.Sones_subtractor.q_RNIIFEO1_3_LC_11_7_4  (
            .in0(N__26223),
            .in1(N__28088),
            .in2(N__26192),
            .in3(N__29812),
            .lcout(\Lab_UT.didp.Sones_subtractor.un8_Mtens_ce ),
            .ltout(\Lab_UT.didp.Sones_subtractor.un8_Mtens_ce_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Sones_subtractor.q_RNIP8IH2_3_LC_11_7_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.Sones_subtractor.q_RNIP8IH2_3_LC_11_7_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Sones_subtractor.q_RNIP8IH2_3_LC_11_7_5 .LUT_INIT=16'b1101111111111111;
    LogicCell40 \Lab_UT.didp.Sones_subtractor.q_RNIP8IH2_3_LC_11_7_5  (
            .in0(N__26795),
            .in1(N__26760),
            .in2(N__26161),
            .in3(N__26678),
            .lcout(\Lab_UT.didp.N_82 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Sones_ce_i_0_o3_LC_11_7_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.Sones_ce_i_0_o3_LC_11_7_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Sones_ce_i_0_o3_LC_11_7_6 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \Lab_UT.didp.Sones_ce_i_0_o3_LC_11_7_6  (
            .in0(N__26679),
            .in1(N__26796),
            .in2(_gnd_net_),
            .in3(N__26761),
            .lcout(\Lab_UT.didp.N_81 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Sones_subtractor.q_RNIVG3M3_3_LC_11_7_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.Sones_subtractor.q_RNIVG3M3_3_LC_11_7_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Sones_subtractor.q_RNIVG3M3_3_LC_11_7_7 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \Lab_UT.didp.Sones_subtractor.q_RNIVG3M3_3_LC_11_7_7  (
            .in0(N__26713),
            .in1(N__26636),
            .in2(N__27091),
            .in3(N__26680),
            .lcout(\Lab_UT.didp.N_83 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Sones_subtractor.q_RNIPVIV3_3_LC_11_8_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.Sones_subtractor.q_RNIPVIV3_3_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Sones_subtractor.q_RNIPVIV3_3_LC_11_8_0 .LUT_INIT=16'b1011111111111111;
    LogicCell40 \Lab_UT.didp.Sones_subtractor.q_RNIPVIV3_3_LC_11_8_0  (
            .in0(N__28049),
            .in1(N__27081),
            .in2(N__28021),
            .in3(N__26638),
            .lcout(\Lab_UT.didp.N_84 ),
            .ltout(\Lab_UT.didp.N_84_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Mtens_subtractor.q_RNI775L5_3_LC_11_8_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mtens_subtractor.q_RNI775L5_3_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Mtens_subtractor.q_RNI775L5_3_LC_11_8_1 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \Lab_UT.didp.Mtens_subtractor.q_RNI775L5_3_LC_11_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26641),
            .in3(N__27046),
            .lcout(\Lab_UT.didp.q_RNI775L5_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Sones_subtractor.q_RNI0E1S4_3_LC_11_8_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.Sones_subtractor.q_RNI0E1S4_3_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Sones_subtractor.q_RNI0E1S4_3_LC_11_8_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.didp.Sones_subtractor.q_RNI0E1S4_3_LC_11_8_2  (
            .in0(N__27044),
            .in1(N__27085),
            .in2(N__28022),
            .in3(N__26637),
            .lcout(\Lab_UT.alarm_match ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Stens_subtractor.q_RNI775L5_3_LC_11_8_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.Stens_subtractor.q_RNI775L5_3_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Stens_subtractor.q_RNI775L5_3_LC_11_8_3 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \Lab_UT.didp.Stens_subtractor.q_RNI775L5_3_LC_11_8_3  (
            .in0(N__28023),
            .in1(N__27043),
            .in2(N__27090),
            .in3(N__28161),
            .lcout(\Lab_UT.didp.Stens_subtractor.q_RNI775L5_0Z0Z_3 ),
            .ltout(\Lab_UT.didp.Stens_subtractor.q_RNI775L5_0Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Stens_subtractor.q_RNO_1_3_LC_11_8_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.Stens_subtractor.q_RNO_1_3_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Stens_subtractor.q_RNO_1_3_LC_11_8_4 .LUT_INIT=16'b0000111100001100;
    LogicCell40 \Lab_UT.didp.Stens_subtractor.q_RNO_1_3_LC_11_8_4  (
            .in0(_gnd_net_),
            .in1(N__27869),
            .in2(N__26605),
            .in3(N__29701),
            .lcout(\Lab_UT.didp.Stens_subtractor.un1_q_c2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Sones_subtractor.q_RNI775L5_3_LC_11_8_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.Sones_subtractor.q_RNI775L5_3_LC_11_8_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Sones_subtractor.q_RNI775L5_3_LC_11_8_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Lab_UT.didp.Sones_subtractor.q_RNI775L5_3_LC_11_8_5  (
            .in0(_gnd_net_),
            .in1(N__28050),
            .in2(_gnd_net_),
            .in3(N__27345),
            .lcout(\Lab_UT.didp.Sones_subtractor.q_RNI775L5_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Stens_subtractor.q_RNO_0_1_LC_11_8_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.Stens_subtractor.q_RNO_0_1_LC_11_8_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Stens_subtractor.q_RNO_0_1_LC_11_8_6 .LUT_INIT=16'b0000010111000101;
    LogicCell40 \Lab_UT.didp.Stens_subtractor.q_RNO_0_1_LC_11_8_6  (
            .in0(N__26583),
            .in1(N__26565),
            .in2(N__28175),
            .in3(N__28818),
            .lcout(\Lab_UT.didp.Stens_subtractor.q_7_i_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Mtens_subtractor.q_RNO_2_1_LC_11_8_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mtens_subtractor.q_RNO_2_1_LC_11_8_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Mtens_subtractor.q_RNO_2_1_LC_11_8_7 .LUT_INIT=16'b1111000011100001;
    LogicCell40 \Lab_UT.didp.Mtens_subtractor.q_RNO_2_1_LC_11_8_7  (
            .in0(N__28684),
            .in1(N__30030),
            .in2(N__27949),
            .in3(N__27045),
            .lcout(\Lab_UT.didp.Mtens_subtractor.q_RNO_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Mtens_subtractor.q_RNO_0_2_LC_11_9_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mtens_subtractor.q_RNO_0_2_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Mtens_subtractor.q_RNO_0_2_LC_11_9_0 .LUT_INIT=16'b1100110010011100;
    LogicCell40 \Lab_UT.didp.Mtens_subtractor.q_RNO_0_2_LC_11_9_0  (
            .in0(N__30028),
            .in1(N__26872),
            .in2(N__26899),
            .in3(N__27943),
            .lcout(),
            .ltout(\Lab_UT.didp.Mtens_subtractor.q_RNO_0_3_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Mtens_subtractor.q_2_LC_11_9_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mtens_subtractor.q_2_LC_11_9_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.Mtens_subtractor.q_2_LC_11_9_1 .LUT_INIT=16'b1111110111101100;
    LogicCell40 \Lab_UT.didp.Mtens_subtractor.q_2_LC_11_9_1  (
            .in0(N__27981),
            .in1(N__26919),
            .in2(N__26974),
            .in3(N__28614),
            .lcout(\Lab_UT.di_Mtens_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29429),
            .ce(),
            .sr(N__28446));
    defparam \Lab_UT.didp.Mtens_subtractor.q_RNIE7IL1_3_LC_11_9_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mtens_subtractor.q_RNIE7IL1_3_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Mtens_subtractor.q_RNIE7IL1_3_LC_11_9_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Lab_UT.didp.Mtens_subtractor.q_RNIE7IL1_3_LC_11_9_2  (
            .in0(N__30027),
            .in1(N__26870),
            .in2(N__26831),
            .in3(N__27942),
            .lcout(\Lab_UT.didp.un3_Mtens_rst ),
            .ltout(\Lab_UT.didp.un3_Mtens_rst_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Mtens_subtractor.q_RNO_0_0_LC_11_9_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mtens_subtractor.q_RNO_0_0_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Mtens_subtractor.q_RNO_0_0_LC_11_9_3 .LUT_INIT=16'b1111110100000010;
    LogicCell40 \Lab_UT.didp.Mtens_subtractor.q_RNO_0_0_LC_11_9_3  (
            .in0(N__28020),
            .in1(N__26961),
            .in2(N__26932),
            .in3(N__30029),
            .lcout(),
            .ltout(\Lab_UT.didp.Mtens_subtractor.un1_q_axb0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Mtens_subtractor.q_0_LC_11_9_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mtens_subtractor.q_0_LC_11_9_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.Mtens_subtractor.q_0_LC_11_9_4 .LUT_INIT=16'b1111101111101010;
    LogicCell40 \Lab_UT.didp.Mtens_subtractor.q_0_LC_11_9_4  (
            .in0(N__26918),
            .in1(N__27980),
            .in2(N__26902),
            .in3(N__29097),
            .lcout(\Lab_UT.didp.di_MtensZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29429),
            .ce(),
            .sr(N__28446));
    defparam \Lab_UT.didp.Stens_subtractor.q_RNI775L5_0_3_LC_11_9_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.Stens_subtractor.q_RNI775L5_0_3_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Stens_subtractor.q_RNI775L5_0_3_LC_11_9_5 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \Lab_UT.didp.Stens_subtractor.q_RNI775L5_0_3_LC_11_9_5  (
            .in0(N__28019),
            .in1(N__27050),
            .in2(N__27089),
            .in3(N__28179),
            .lcout(\Lab_UT.didp.Mtens_ce ),
            .ltout(\Lab_UT.didp.Mtens_ce_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Mtens_subtractor.q_RNO_0_3_LC_11_9_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mtens_subtractor.q_RNO_0_3_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Mtens_subtractor.q_RNO_0_3_LC_11_9_6 .LUT_INIT=16'b1010011010011010;
    LogicCell40 \Lab_UT.didp.Mtens_subtractor.q_RNO_0_3_LC_11_9_6  (
            .in0(N__26824),
            .in1(N__26871),
            .in2(N__26839),
            .in3(N__27958),
            .lcout(),
            .ltout(\Lab_UT.didp.Mtens_subtractor.q_RNO_0_2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Mtens_subtractor.q_3_LC_11_9_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mtens_subtractor.q_3_LC_11_9_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.Mtens_subtractor.q_3_LC_11_9_7 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \Lab_UT.didp.Mtens_subtractor.q_3_LC_11_9_7  (
            .in0(N__27982),
            .in1(_gnd_net_),
            .in2(N__26836),
            .in3(N__28987),
            .lcout(\Lab_UT.didp.di_Mtens_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29429),
            .ce(),
            .sr(N__28446));
    defparam \Lab_UT.didp.Mones_subtractor.q_RNIN8C59_3_LC_11_10_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mones_subtractor.q_RNIN8C59_3_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Mones_subtractor.q_RNIN8C59_3_LC_11_10_0 .LUT_INIT=16'b1100010010000000;
    LogicCell40 \Lab_UT.didp.Mones_subtractor.q_RNIN8C59_3_LC_11_10_0  (
            .in0(N__29950),
            .in1(N__30107),
            .in2(N__27325),
            .in3(N__27435),
            .lcout(\Lab_UT.didp.Mones_subtractor.q_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.dicLdMones_LC_11_10_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.dicLdMones_LC_11_10_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.dicLdMones_LC_11_10_1 .LUT_INIT=16'b1100101011001100;
    LogicCell40 \Lab_UT.dictrl.dicLdMones_LC_11_10_1  (
            .in0(N__27436),
            .in1(N__27324),
            .in2(N__29962),
            .in3(N__29891),
            .lcout(\Lab_UT.dicLdMones ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29420),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.dicLdMtens_LC_11_10_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.dicLdMtens_LC_11_10_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.dicLdMtens_LC_11_10_2 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \Lab_UT.dictrl.dicLdMtens_LC_11_10_2  (
            .in0(N__29892),
            .in1(N__27006),
            .in2(N__26992),
            .in3(N__29956),
            .lcout(\Lab_UT.dicLdMtens ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29420),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_0_ret_6_RNIU5JA3_LC_11_10_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_6_RNIU5JA3_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_0_ret_6_RNIU5JA3_LC_11_10_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_6_RNIU5JA3_LC_11_10_3  (
            .in0(N__27313),
            .in1(N__27813),
            .in2(_gnd_net_),
            .in3(N__27301),
            .lcout(\Lab_UT.dicLdMtens_latmux ),
            .ltout(\Lab_UT.dicLdMtens_latmux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Mtens_subtractor.q_7_i_o2_2_LC_11_10_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mtens_subtractor.q_7_i_o2_2_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Mtens_subtractor.q_7_i_o2_2_LC_11_10_4 .LUT_INIT=16'b0010011111111111;
    LogicCell40 \Lab_UT.didp.Mtens_subtractor.q_7_i_o2_2_LC_11_10_4  (
            .in0(N__29951),
            .in1(N__27002),
            .in2(N__27169),
            .in3(N__28682),
            .lcout(\Lab_UT.didp.Mtens_subtractor.N_87 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Stens_subtractor.q_RNI68H41_3_LC_11_10_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.Stens_subtractor.q_RNI68H41_3_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Stens_subtractor.q_RNI68H41_3_LC_11_10_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Lab_UT.didp.Stens_subtractor.q_RNI68H41_3_LC_11_10_5  (
            .in0(N__27166),
            .in1(N__27870),
            .in2(N__27130),
            .in3(N__29699),
            .lcout(\Lab_UT.didp.un6_Mtens_ce ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Mtens_subtractor.q_RNO_0_1_LC_11_10_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mtens_subtractor.q_RNO_0_1_LC_11_10_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Mtens_subtractor.q_RNO_0_1_LC_11_10_6 .LUT_INIT=16'b0000000010111110;
    LogicCell40 \Lab_UT.didp.Mtens_subtractor.q_RNO_0_1_LC_11_10_6  (
            .in0(N__27051),
            .in1(N__30037),
            .in2(N__27947),
            .in3(N__28683),
            .lcout(\Lab_UT.didp.Mtens_subtractor.N_145 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Mtens_subtractor.q_RNO_1_1_LC_11_10_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mtens_subtractor.q_RNO_1_1_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Mtens_subtractor.q_RNO_1_1_LC_11_10_7 .LUT_INIT=16'b0000001000010011;
    LogicCell40 \Lab_UT.didp.Mtens_subtractor.q_RNO_1_1_LC_11_10_7  (
            .in0(N__29952),
            .in1(N__27016),
            .in2(N__27007),
            .in3(N__26988),
            .lcout(\Lab_UT.didp.Mtens_subtractor.N_147 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Mtens_subtractor.q_1_LC_11_11_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mtens_subtractor.q_1_LC_11_11_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.Mtens_subtractor.q_1_LC_11_11_0 .LUT_INIT=16'b0000000001010100;
    LogicCell40 \Lab_UT.didp.Mtens_subtractor.q_1_LC_11_11_0  (
            .in0(N__26980),
            .in1(N__27979),
            .in2(N__28822),
            .in3(N__27964),
            .lcout(\Lab_UT.didp.di_Mtens_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29412),
            .ce(),
            .sr(N__28456));
    defparam \Lab_UT.didp.Mtens_subtractor.q_RNO_1_3_LC_11_11_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mtens_subtractor.q_RNO_1_3_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Mtens_subtractor.q_RNO_1_3_LC_11_11_1 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \Lab_UT.didp.Mtens_subtractor.q_RNO_1_3_LC_11_11_1  (
            .in0(N__28678),
            .in1(N__30039),
            .in2(_gnd_net_),
            .in3(N__27934),
            .lcout(\Lab_UT.didp.Mtens_subtractor.un1_q_c2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Mones_subtractor.q_RNITOVP_1_LC_11_11_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mones_subtractor.q_RNITOVP_1_LC_11_11_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Mones_subtractor.q_RNITOVP_1_LC_11_11_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \Lab_UT.didp.Mones_subtractor.q_RNITOVP_1_LC_11_11_2  (
            .in0(N__30081),
            .in1(N__27938),
            .in2(_gnd_net_),
            .in3(N__29780),
            .lcout(),
            .ltout(\Lab_UT.didp.q_RNITOVP_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.curr_LED_RNIJFM52_1_LC_11_11_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.curr_LED_RNIJFM52_1_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.curr_LED_RNIJFM52_1_LC_11_11_3 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \Lab_UT.didp.curr_LED_RNIJFM52_1_LC_11_11_3  (
            .in0(N__27832),
            .in1(_gnd_net_),
            .in2(N__27892),
            .in3(N__29644),
            .lcout(led_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Stens_subtractor.q_RNI99F11_1_LC_11_11_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.Stens_subtractor.q_RNI99F11_1_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Stens_subtractor.q_RNI99F11_1_LC_11_11_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Lab_UT.didp.Stens_subtractor.q_RNI99F11_1_LC_11_11_4  (
            .in0(N__27871),
            .in1(N__29781),
            .in2(_gnd_net_),
            .in3(N__28105),
            .lcout(\Lab_UT.didp.q_RNI99F11_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.currState_0_ret_12_RNIB2D93_LC_11_12_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.currState_0_ret_12_RNIB2D93_LC_11_12_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.currState_0_ret_12_RNIB2D93_LC_11_12_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.dictrl.currState_0_ret_12_RNIB2D93_LC_11_12_3  (
            .in0(N__27826),
            .in1(N__27812),
            .in2(_gnd_net_),
            .in3(N__27562),
            .lcout(\Lab_UT.dicLdMones_latmux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.displayAlarm_6_LC_12_4_0 .C_ON=1'b0;
    defparam \Lab_UT.displayAlarm_6_LC_12_4_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.displayAlarm_6_LC_12_4_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Lab_UT.displayAlarm_6_LC_12_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29532),
            .lcout(\Lab_UT.displayAlarmZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29474),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.displayAlarm_4_LC_12_5_1 .C_ON=1'b0;
    defparam \Lab_UT.displayAlarm_4_LC_12_5_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.displayAlarm_4_LC_12_5_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Lab_UT.displayAlarm_4_LC_12_5_1  (
            .in0(_gnd_net_),
            .in1(N__29546),
            .in2(_gnd_net_),
            .in3(N__27413),
            .lcout(\Lab_UT.displayAlarmZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29467),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Sones_subtractor.q_RNO_1_1_LC_12_7_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.Sones_subtractor.q_RNO_1_1_LC_12_7_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Sones_subtractor.q_RNO_1_1_LC_12_7_0 .LUT_INIT=16'b1100110011001001;
    LogicCell40 \Lab_UT.didp.Sones_subtractor.q_RNO_1_1_LC_12_7_0  (
            .in0(N__27341),
            .in1(N__28092),
            .in2(N__28059),
            .in3(N__29814),
            .lcout(\Lab_UT.didp.Sones_subtractor.q_RNO_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.dicLdSones_RNISPBP3_LC_12_7_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.dicLdSones_RNISPBP3_LC_12_7_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.dicLdSones_RNISPBP3_LC_12_7_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \Lab_UT.dictrl.dicLdSones_RNISPBP3_LC_12_7_1  (
            .in0(N__29961),
            .in1(_gnd_net_),
            .in2(N__29845),
            .in3(N__29867),
            .lcout(),
            .ltout(\Lab_UT.ld_enable_Sones_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Sones_subtractor.q_RNO_0_1_LC_12_7_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.Sones_subtractor.q_RNO_0_1_LC_12_7_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Sones_subtractor.q_RNO_0_1_LC_12_7_2 .LUT_INIT=16'b0000000001011111;
    LogicCell40 \Lab_UT.didp.Sones_subtractor.q_RNO_0_1_LC_12_7_2  (
            .in0(N__28055),
            .in1(_gnd_net_),
            .in2(N__28210),
            .in3(N__28207),
            .lcout(),
            .ltout(\Lab_UT.didp.Sones_subtractor.q_7_i_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Sones_subtractor.q_1_LC_12_7_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.Sones_subtractor.q_1_LC_12_7_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.Sones_subtractor.q_1_LC_12_7_3 .LUT_INIT=16'b0000110000001000;
    LogicCell40 \Lab_UT.didp.Sones_subtractor.q_1_LC_12_7_3  (
            .in0(N__28124),
            .in1(N__28174),
            .in2(N__28201),
            .in3(N__28820),
            .lcout(\Lab_UT.didp.di_Sones_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29452),
            .ce(),
            .sr(N__28455));
    defparam \Lab_UT.didp.Sones_subtractor.q_RNO_0_0_LC_12_7_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.Sones_subtractor.q_RNO_0_0_LC_12_7_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Sones_subtractor.q_RNO_0_0_LC_12_7_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \Lab_UT.didp.Sones_subtractor.q_RNO_0_0_LC_12_7_4  (
            .in0(_gnd_net_),
            .in1(N__28198),
            .in2(_gnd_net_),
            .in3(N__29816),
            .lcout(),
            .ltout(\Lab_UT.didp.Sones_subtractor.un1_q_axb0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Sones_subtractor.q_0_LC_12_7_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.Sones_subtractor.q_0_LC_12_7_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.Sones_subtractor.q_0_LC_12_7_5 .LUT_INIT=16'b1111011110110011;
    LogicCell40 \Lab_UT.didp.Sones_subtractor.q_0_LC_12_7_5  (
            .in0(N__28123),
            .in1(N__28173),
            .in2(N__28129),
            .in3(N__29107),
            .lcout(\Lab_UT.didp.di_Sones_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29452),
            .ce(),
            .sr(N__28455));
    defparam \Lab_UT.didp.Sones_subtractor.q_7_i_o2_3_LC_12_7_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.Sones_subtractor.q_7_i_o2_3_LC_12_7_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Sones_subtractor.q_7_i_o2_3_LC_12_7_6 .LUT_INIT=16'b0011111101011111;
    LogicCell40 \Lab_UT.didp.Sones_subtractor.q_7_i_o2_3_LC_12_7_6  (
            .in0(N__29868),
            .in1(N__29843),
            .in2(N__28060),
            .in3(N__29960),
            .lcout(\Lab_UT.didp.Sones_subtractor.N_85 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Sones_subtractor.q_RNO_1_3_LC_12_7_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.Sones_subtractor.q_RNO_1_3_LC_12_7_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Sones_subtractor.q_RNO_1_3_LC_12_7_7 .LUT_INIT=16'b0000000011111010;
    LogicCell40 \Lab_UT.didp.Sones_subtractor.q_RNO_1_3_LC_12_7_7  (
            .in0(N__29815),
            .in1(_gnd_net_),
            .in2(N__28103),
            .in3(N__28051),
            .lcout(\Lab_UT.didp.Sones_subtractor.un1_q_c2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Mones_subtractor.q_RNIQEF9_3_LC_12_8_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mones_subtractor.q_RNIQEF9_3_LC_12_8_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Mones_subtractor.q_RNIQEF9_3_LC_12_8_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Lab_UT.didp.Mones_subtractor.q_RNIQEF9_3_LC_12_8_0  (
            .in0(N__28285),
            .in1(N__30072),
            .in2(N__28247),
            .in3(N__29985),
            .lcout(\Lab_UT.didp.un4_Mtens_ce ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Mones_subtractor.q_RNO_0_0_LC_12_8_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mones_subtractor.q_RNO_0_0_LC_12_8_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Mones_subtractor.q_RNO_0_0_LC_12_8_1 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \Lab_UT.didp.Mones_subtractor.q_RNO_0_0_LC_12_8_1  (
            .in0(N__29986),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30120),
            .lcout(),
            .ltout(\Lab_UT.didp.Mones_subtractor.un1_q_axb_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Mones_subtractor.q_0_LC_12_8_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mones_subtractor.q_0_LC_12_8_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.Mones_subtractor.q_0_LC_12_8_2 .LUT_INIT=16'b1111110101110101;
    LogicCell40 \Lab_UT.didp.Mones_subtractor.q_0_LC_12_8_2  (
            .in0(N__28660),
            .in1(N__28633),
            .in2(N__29110),
            .in3(N__29098),
            .lcout(\Lab_UT.didp.di_Mones_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29444),
            .ce(),
            .sr(N__28447));
    defparam \Lab_UT.didp.Mones_subtractor.q_3_LC_12_8_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mones_subtractor.q_3_LC_12_8_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.Mones_subtractor.q_3_LC_12_8_3 .LUT_INIT=16'b1111101101110011;
    LogicCell40 \Lab_UT.didp.Mones_subtractor.q_3_LC_12_8_3  (
            .in0(N__28636),
            .in1(N__28665),
            .in2(N__30136),
            .in3(N__28980),
            .lcout(\Lab_UT.didp.di_Mones_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29444),
            .ce(),
            .sr(N__28447));
    defparam \Lab_UT.didp.Mones_subtractor.q_1_LC_12_8_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mones_subtractor.q_1_LC_12_8_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.Mones_subtractor.q_1_LC_12_8_4 .LUT_INIT=16'b1110000000100000;
    LogicCell40 \Lab_UT.didp.Mones_subtractor.q_1_LC_12_8_4  (
            .in0(N__30046),
            .in1(N__28634),
            .in2(N__28677),
            .in3(N__28819),
            .lcout(\Lab_UT.didp.di_Mones_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29444),
            .ce(),
            .sr(N__28447));
    defparam \Lab_UT.didp.Mones_subtractor.q_RNO_0_2_LC_12_8_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mones_subtractor.q_RNO_0_2_LC_12_8_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Mones_subtractor.q_RNO_0_2_LC_12_8_5 .LUT_INIT=16'b1110111000010001;
    LogicCell40 \Lab_UT.didp.Mones_subtractor.q_RNO_0_2_LC_12_8_5  (
            .in0(N__28264),
            .in1(N__30121),
            .in2(_gnd_net_),
            .in3(N__28286),
            .lcout(),
            .ltout(\Lab_UT.didp.Mones_subtractor.q_RNO_0_2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Mones_subtractor.q_2_LC_12_8_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mones_subtractor.q_2_LC_12_8_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.Mones_subtractor.q_2_LC_12_8_6 .LUT_INIT=16'b1010100000100000;
    LogicCell40 \Lab_UT.didp.Mones_subtractor.q_2_LC_12_8_6  (
            .in0(N__28664),
            .in1(N__28635),
            .in2(N__28618),
            .in3(N__28607),
            .lcout(\Lab_UT.didp.di_Mones_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29444),
            .ce(),
            .sr(N__28447));
    defparam \Lab_UT.didp.Mones_subtractor.un1_q_cry_0_s1_c_LC_12_9_0 .C_ON=1'b1;
    defparam \Lab_UT.didp.Mones_subtractor.un1_q_cry_0_s1_c_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Mones_subtractor.un1_q_cry_0_s1_c_LC_12_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \Lab_UT.didp.Mones_subtractor.un1_q_cry_0_s1_c_LC_12_9_0  (
            .in0(_gnd_net_),
            .in1(N__29987),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_9_0_),
            .carryout(\Lab_UT.didp.Mones_subtractor.un1_q_cry_0_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Mones_subtractor.un1_q_cry_0_s1_THRU_LUT4_0_LC_12_9_1 .C_ON=1'b1;
    defparam \Lab_UT.didp.Mones_subtractor.un1_q_cry_0_s1_THRU_LUT4_0_LC_12_9_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Mones_subtractor.un1_q_cry_0_s1_THRU_LUT4_0_LC_12_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.Mones_subtractor.un1_q_cry_0_s1_THRU_LUT4_0_LC_12_9_1  (
            .in0(_gnd_net_),
            .in1(N__30073),
            .in2(N__28357),
            .in3(N__28360),
            .lcout(\Lab_UT.didp.Mones_subtractor.un1_q_cry_0_s1_THRU_CO ),
            .ltout(),
            .carryin(\Lab_UT.didp.Mones_subtractor.un1_q_cry_0_s1 ),
            .carryout(\Lab_UT.didp.Mones_subtractor.un1_q_cry_1_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Mones_subtractor.un1_q_cry_1_s1_THRU_LUT4_0_LC_12_9_2 .C_ON=1'b1;
    defparam \Lab_UT.didp.Mones_subtractor.un1_q_cry_1_s1_THRU_LUT4_0_LC_12_9_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Mones_subtractor.un1_q_cry_1_s1_THRU_LUT4_0_LC_12_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.Mones_subtractor.un1_q_cry_1_s1_THRU_LUT4_0_LC_12_9_2  (
            .in0(_gnd_net_),
            .in1(N__28353),
            .in2(N__28295),
            .in3(N__28255),
            .lcout(\Lab_UT.didp.Mones_subtractor.un1_q_cry_1_s1_THRU_CO ),
            .ltout(),
            .carryin(\Lab_UT.didp.Mones_subtractor.un1_q_cry_1_s1 ),
            .carryout(\Lab_UT.didp.Mones_subtractor.un1_q_cry_2_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Mones_subtractor.q_RNO_0_3_LC_12_9_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mones_subtractor.q_RNO_0_3_LC_12_9_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Mones_subtractor.q_RNO_0_3_LC_12_9_3 .LUT_INIT=16'b1010101010011001;
    LogicCell40 \Lab_UT.didp.Mones_subtractor.q_RNO_0_3_LC_12_9_3  (
            .in0(N__28240),
            .in1(N__30119),
            .in2(_gnd_net_),
            .in3(N__28213),
            .lcout(\Lab_UT.didp.Mones_subtractor.q_RNO_0_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Mones_subtractor.q_RNO_0_1_LC_12_9_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mones_subtractor.q_RNO_0_1_LC_12_9_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Mones_subtractor.q_RNO_0_1_LC_12_9_5 .LUT_INIT=16'b1110111000010001;
    LogicCell40 \Lab_UT.didp.Mones_subtractor.q_RNO_0_1_LC_12_9_5  (
            .in0(N__30127),
            .in1(N__30118),
            .in2(_gnd_net_),
            .in3(N__30074),
            .lcout(\Lab_UT.didp.Mones_subtractor.q_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Mones_subtractor.q_RNIRMVP_0_LC_12_9_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.Mones_subtractor.q_RNIRMVP_0_LC_12_9_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Mones_subtractor.q_RNIRMVP_0_LC_12_9_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Lab_UT.didp.Mones_subtractor.q_RNIRMVP_0_LC_12_9_6  (
            .in0(N__30040),
            .in1(N__29774),
            .in2(_gnd_net_),
            .in3(N__29988),
            .lcout(\Lab_UT.didp.q_RNIRMVP_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.dicLdSones_LC_12_10_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.dicLdSones_LC_12_10_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.dicLdSones_LC_12_10_4 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \Lab_UT.dictrl.dicLdSones_LC_12_10_4  (
            .in0(N__29957),
            .in1(N__29893),
            .in2(N__29844),
            .in3(N__29869),
            .lcout(\Lab_UT.dicLdSones ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29430),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.Stens_subtractor.q_RNI77F11_0_LC_12_10_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.Stens_subtractor.q_RNI77F11_0_LC_12_10_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.Stens_subtractor.q_RNI77F11_0_LC_12_10_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \Lab_UT.didp.Stens_subtractor.q_RNI77F11_0_LC_12_10_6  (
            .in0(N__29821),
            .in1(N__29782),
            .in2(_gnd_net_),
            .in3(N__29700),
            .lcout(),
            .ltout(\Lab_UT.didp.q_RNI77F11_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.curr_LED_RNIFBM52_1_LC_12_10_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.curr_LED_RNIFBM52_1_LC_12_10_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.curr_LED_RNIFBM52_1_LC_12_10_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \Lab_UT.didp.curr_LED_RNIFBM52_1_LC_12_10_7  (
            .in0(_gnd_net_),
            .in1(N__29653),
            .in2(N__29647),
            .in3(N__29637),
            .lcout(led_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.r_dicAlarmIdle_LC_12_11_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.r_dicAlarmIdle_LC_12_11_0 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.r_dicAlarmIdle_LC_12_11_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.dictrl.r_dicAlarmIdle_LC_12_11_0  (
            .in0(_gnd_net_),
            .in1(N__29512),
            .in2(_gnd_net_),
            .in3(N__29584),
            .lcout(\Lab_UT.alarm_off ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__29421),
            .ce(),
            .sr(N__29131));
endmodule // latticehx1k
